// soc_system.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module soc_system (
		output wire [2:0]  button_pio_external_connection_export,  // button_pio_external_connection.export
		input  wire        clk_50_clk,                             //                         clk_50.clk
		input  wire        clk_cnn_clk,                            //                        clk_cnn.clk
		output wire [2:0]  dipsw_pio_external_connection_export,   //  dipsw_pio_external_connection.export
		input  wire        hps_0_f2h_cold_reset_req_reset_n,       //       hps_0_f2h_cold_reset_req.reset_n
		input  wire        hps_0_f2h_debug_reset_req_reset_n,      //      hps_0_f2h_debug_reset_req.reset_n
		input  wire [27:0] hps_0_f2h_stm_hw_events_stm_hwevents,   //        hps_0_f2h_stm_hw_events.stm_hwevents
		input  wire        hps_0_f2h_warm_reset_req_reset_n,       //       hps_0_f2h_warm_reset_req.reset_n
		output wire [66:0] hps_0_h2f_loan_io_in,                   //              hps_0_h2f_loan_io.in
		input  wire [66:0] hps_0_h2f_loan_io_out,                  //                               .out
		input  wire [66:0] hps_0_h2f_loan_io_oe,                   //                               .oe
		output wire        hps_0_h2f_reset_reset_n,                //                hps_0_h2f_reset.reset_n
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CLK,  //                   hps_0_hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD0,    //                               .hps_io_emac1_inst_TXD0
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD1,    //                               .hps_io_emac1_inst_TXD1
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD2,    //                               .hps_io_emac1_inst_TXD2
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD3,    //                               .hps_io_emac1_inst_TXD3
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD0,    //                               .hps_io_emac1_inst_RXD0
		inout  wire        hps_0_hps_io_hps_io_emac1_inst_MDIO,    //                               .hps_io_emac1_inst_MDIO
		output wire        hps_0_hps_io_hps_io_emac1_inst_MDC,     //                               .hps_io_emac1_inst_MDC
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CTL,  //                               .hps_io_emac1_inst_RX_CTL
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CTL,  //                               .hps_io_emac1_inst_TX_CTL
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CLK,  //                               .hps_io_emac1_inst_RX_CLK
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD1,    //                               .hps_io_emac1_inst_RXD1
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD2,    //                               .hps_io_emac1_inst_RXD2
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD3,    //                               .hps_io_emac1_inst_RXD3
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_CMD,      //                               .hps_io_sdio_inst_CMD
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D0,       //                               .hps_io_sdio_inst_D0
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D1,       //                               .hps_io_sdio_inst_D1
		output wire        hps_0_hps_io_hps_io_sdio_inst_CLK,      //                               .hps_io_sdio_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D2,       //                               .hps_io_sdio_inst_D2
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D3,       //                               .hps_io_sdio_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D0,       //                               .hps_io_usb1_inst_D0
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D1,       //                               .hps_io_usb1_inst_D1
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D2,       //                               .hps_io_usb1_inst_D2
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D3,       //                               .hps_io_usb1_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D4,       //                               .hps_io_usb1_inst_D4
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D5,       //                               .hps_io_usb1_inst_D5
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D6,       //                               .hps_io_usb1_inst_D6
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D7,       //                               .hps_io_usb1_inst_D7
		input  wire        hps_0_hps_io_hps_io_usb1_inst_CLK,      //                               .hps_io_usb1_inst_CLK
		output wire        hps_0_hps_io_hps_io_usb1_inst_STP,      //                               .hps_io_usb1_inst_STP
		input  wire        hps_0_hps_io_hps_io_usb1_inst_DIR,      //                               .hps_io_usb1_inst_DIR
		input  wire        hps_0_hps_io_hps_io_usb1_inst_NXT,      //                               .hps_io_usb1_inst_NXT
		input  wire        hps_0_hps_io_hps_io_uart0_inst_RX,      //                               .hps_io_uart0_inst_RX
		output wire        hps_0_hps_io_hps_io_uart0_inst_TX,      //                               .hps_io_uart0_inst_TX
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO34,   //                               .hps_io_gpio_inst_GPIO34
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO35,   //                               .hps_io_gpio_inst_GPIO35
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO48,   //                               .hps_io_gpio_inst_GPIO48
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO51,   //                               .hps_io_gpio_inst_GPIO51
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO52,   //                               .hps_io_gpio_inst_GPIO52
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO53,   //                               .hps_io_gpio_inst_GPIO53
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO54,   //                               .hps_io_gpio_inst_GPIO54
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_LOANIO00, //                               .hps_io_gpio_inst_LOANIO00
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_LOANIO09, //                               .hps_io_gpio_inst_LOANIO09
		input  wire [19:0] led_pio_external_connection_export,     //    led_pio_external_connection.export
		output wire [14:0] memory_mem_a,                           //                         memory.mem_a
		output wire [2:0]  memory_mem_ba,                          //                               .mem_ba
		output wire        memory_mem_ck,                          //                               .mem_ck
		output wire        memory_mem_ck_n,                        //                               .mem_ck_n
		output wire        memory_mem_cke,                         //                               .mem_cke
		output wire        memory_mem_cs_n,                        //                               .mem_cs_n
		output wire        memory_mem_ras_n,                       //                               .mem_ras_n
		output wire        memory_mem_cas_n,                       //                               .mem_cas_n
		output wire        memory_mem_we_n,                        //                               .mem_we_n
		output wire        memory_mem_reset_n,                     //                               .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                          //                               .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                         //                               .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                       //                               .mem_dqs_n
		output wire        memory_mem_odt,                         //                               .mem_odt
		output wire [3:0]  memory_mem_dm,                          //                               .mem_dm
		input  wire        memory_oct_rzqin,                       //                               .oct_rzqin
		input  wire        reset_50_reset_n,                       //                       reset_50.reset_n
		input  wire        reset_cnn_reset_n                       //                      reset_cnn.reset_n
	);

	wire          vcam_0_dvp_bus_dvp_pclk;                                        // vcam_0:dvp_pclk -> dvp_ddr3_0:dvp_pclk
	wire          vcam_0_dvp_bus_dvp_vsync;                                       // vcam_0:dvp_vsync -> dvp_ddr3_0:dvp_vsync
	wire          vcam_0_dvp_bus_dvp_href;                                        // vcam_0:dvp_href -> dvp_ddr3_0:dvp_href
	wire    [7:0] vcam_0_dvp_bus_dvp_data;                                        // vcam_0:dvp_data -> dvp_ddr3_0:dvp_data
	wire          ddr3_vga_0_vga_bus_vga_vsync;                                   // ddr3_vga_0:vga_vsync -> vhdmi_0:vga_vsync
	wire          ddr3_vga_0_vga_bus_vga_de;                                      // ddr3_vga_0:vga_de -> vhdmi_0:vga_de
	wire          ddr3_vga_0_vga_bus_vga_clk;                                     // ddr3_vga_0:vga_clk -> vhdmi_0:vga_clk
	wire          ddr3_vga_0_vga_bus_vga_hsync;                                   // ddr3_vga_0:vga_hsync -> vhdmi_0:vga_hsync
	wire   [23:0] ddr3_vga_0_vga_bus_vga_rgb;                                     // ddr3_vga_0:vga_rgb -> vhdmi_0:vga_rgb
	wire          vcam_0_data_bus_waitrequest;                                    // mm_interconnect_0:vcam_0_data_bus_waitrequest -> vcam_0:avm_waitrequest
	wire  [127:0] vcam_0_data_bus_readdata;                                       // mm_interconnect_0:vcam_0_data_bus_readdata -> vcam_0:avm_rdata
	wire          vcam_0_data_bus_read;                                           // vcam_0:avm_read -> mm_interconnect_0:vcam_0_data_bus_read
	wire   [31:0] vcam_0_data_bus_address;                                        // vcam_0:avm_addr -> mm_interconnect_0:vcam_0_data_bus_address
	wire   [15:0] vcam_0_data_bus_byteenable;                                     // vcam_0:avm_byteenable -> mm_interconnect_0:vcam_0_data_bus_byteenable
	wire          vcam_0_data_bus_readdatavalid;                                  // mm_interconnect_0:vcam_0_data_bus_readdatavalid -> vcam_0:avm_rdata_valid
	wire          vcam_0_data_bus_write;                                          // vcam_0:avm_write -> mm_interconnect_0:vcam_0_data_bus_write
	wire  [127:0] vcam_0_data_bus_writedata;                                      // vcam_0:avm_wdata -> mm_interconnect_0:vcam_0_data_bus_writedata
	wire    [9:0] vcam_0_data_bus_burstcount;                                     // vcam_0:avm_size -> mm_interconnect_0:vcam_0_data_bus_burstcount
	wire          dvp_ddr3_0_data_bus_waitrequest;                                // mm_interconnect_0:dvp_ddr3_0_data_bus_waitrequest -> dvp_ddr3_0:avl_waitrequest
	wire  [127:0] dvp_ddr3_0_data_bus_readdata;                                   // mm_interconnect_0:dvp_ddr3_0_data_bus_readdata -> dvp_ddr3_0:avl_rdata
	wire   [31:0] dvp_ddr3_0_data_bus_address;                                    // dvp_ddr3_0:avl_addr -> mm_interconnect_0:dvp_ddr3_0_data_bus_address
	wire   [15:0] dvp_ddr3_0_data_bus_byteenable;                                 // dvp_ddr3_0:avl_be -> mm_interconnect_0:dvp_ddr3_0_data_bus_byteenable
	wire          dvp_ddr3_0_data_bus_read;                                       // dvp_ddr3_0:avl_read_req -> mm_interconnect_0:dvp_ddr3_0_data_bus_read
	wire          dvp_ddr3_0_data_bus_readdatavalid;                              // mm_interconnect_0:dvp_ddr3_0_data_bus_readdatavalid -> dvp_ddr3_0:avl_rdata_valid
	wire  [127:0] dvp_ddr3_0_data_bus_writedata;                                  // dvp_ddr3_0:avl_wdata -> mm_interconnect_0:dvp_ddr3_0_data_bus_writedata
	wire          dvp_ddr3_0_data_bus_write;                                      // dvp_ddr3_0:avl_write_req -> mm_interconnect_0:dvp_ddr3_0_data_bus_write
	wire    [9:0] dvp_ddr3_0_data_bus_burstcount;                                 // dvp_ddr3_0:avl_size -> mm_interconnect_0:dvp_ddr3_0_data_bus_burstcount
	wire          ddr3_vga_0_data_bus_waitrequest;                                // mm_interconnect_0:ddr3_vga_0_data_bus_waitrequest -> ddr3_vga_0:avl_waitrequest
	wire  [127:0] ddr3_vga_0_data_bus_readdata;                                   // mm_interconnect_0:ddr3_vga_0_data_bus_readdata -> ddr3_vga_0:avl_rdata
	wire   [31:0] ddr3_vga_0_data_bus_address;                                    // ddr3_vga_0:avl_addr -> mm_interconnect_0:ddr3_vga_0_data_bus_address
	wire   [15:0] ddr3_vga_0_data_bus_byteenable;                                 // ddr3_vga_0:avl_be -> mm_interconnect_0:ddr3_vga_0_data_bus_byteenable
	wire          ddr3_vga_0_data_bus_read;                                       // ddr3_vga_0:avl_read_req -> mm_interconnect_0:ddr3_vga_0_data_bus_read
	wire          ddr3_vga_0_data_bus_readdatavalid;                              // mm_interconnect_0:ddr3_vga_0_data_bus_readdatavalid -> ddr3_vga_0:avl_rdata_valid
	wire  [127:0] ddr3_vga_0_data_bus_writedata;                                  // ddr3_vga_0:avl_wdata -> mm_interconnect_0:ddr3_vga_0_data_bus_writedata
	wire          ddr3_vga_0_data_bus_write;                                      // ddr3_vga_0:avl_write_req -> mm_interconnect_0:ddr3_vga_0_data_bus_write
	wire    [9:0] ddr3_vga_0_data_bus_burstcount;                                 // ddr3_vga_0:avl_size -> mm_interconnect_0:ddr3_vga_0_data_bus_burstcount
	wire          vhdmi_0_m_avalon_mm_waitrequest;                                // mm_interconnect_0:vhdmi_0_m_avalon_mm_waitrequest -> vhdmi_0:m_avl_waitrequest
	wire   [31:0] vhdmi_0_m_avalon_mm_address;                                    // vhdmi_0:m_avl_addr -> mm_interconnect_0:vhdmi_0_m_avalon_mm_address
	wire   [15:0] vhdmi_0_m_avalon_mm_byteenable;                                 // vhdmi_0:m_avl_be -> mm_interconnect_0:vhdmi_0_m_avalon_mm_byteenable
	wire  [127:0] vhdmi_0_m_avalon_mm_writedata;                                  // vhdmi_0:m_avl_wdata -> mm_interconnect_0:vhdmi_0_m_avalon_mm_writedata
	wire          vhdmi_0_m_avalon_mm_write;                                      // vhdmi_0:m_avl_write_req -> mm_interconnect_0:vhdmi_0_m_avalon_mm_write
	wire    [7:0] vhdmi_0_m_avalon_mm_burstcount;                                 // vhdmi_0:m_avl_size -> mm_interconnect_0:vhdmi_0_m_avalon_mm_burstcount
	wire  [127:0] mm_interconnect_0_mm_bridge_axi_s0_readdata;                    // mm_bridge_axi:s0_readdata -> mm_interconnect_0:mm_bridge_axi_s0_readdata
	wire          mm_interconnect_0_mm_bridge_axi_s0_waitrequest;                 // mm_bridge_axi:s0_waitrequest -> mm_interconnect_0:mm_bridge_axi_s0_waitrequest
	wire          mm_interconnect_0_mm_bridge_axi_s0_debugaccess;                 // mm_interconnect_0:mm_bridge_axi_s0_debugaccess -> mm_bridge_axi:s0_debugaccess
	wire   [31:0] mm_interconnect_0_mm_bridge_axi_s0_address;                     // mm_interconnect_0:mm_bridge_axi_s0_address -> mm_bridge_axi:s0_address
	wire          mm_interconnect_0_mm_bridge_axi_s0_read;                        // mm_interconnect_0:mm_bridge_axi_s0_read -> mm_bridge_axi:s0_read
	wire   [15:0] mm_interconnect_0_mm_bridge_axi_s0_byteenable;                  // mm_interconnect_0:mm_bridge_axi_s0_byteenable -> mm_bridge_axi:s0_byteenable
	wire          mm_interconnect_0_mm_bridge_axi_s0_readdatavalid;               // mm_bridge_axi:s0_readdatavalid -> mm_interconnect_0:mm_bridge_axi_s0_readdatavalid
	wire          mm_interconnect_0_mm_bridge_axi_s0_write;                       // mm_interconnect_0:mm_bridge_axi_s0_write -> mm_bridge_axi:s0_write
	wire  [127:0] mm_interconnect_0_mm_bridge_axi_s0_writedata;                   // mm_interconnect_0:mm_bridge_axi_s0_writedata -> mm_bridge_axi:s0_writedata
	wire    [4:0] mm_interconnect_0_mm_bridge_axi_s0_burstcount;                  // mm_interconnect_0:mm_bridge_axi_s0_burstcount -> mm_bridge_axi:s0_burstcount
	wire    [1:0] hps_0_h2f_lw_axi_master_awburst;                                // hps_0:h2f_lw_AWBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awburst
	wire    [3:0] hps_0_h2f_lw_axi_master_arlen;                                  // hps_0:h2f_lw_ARLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlen
	wire    [3:0] hps_0_h2f_lw_axi_master_wstrb;                                  // hps_0:h2f_lw_WSTRB -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wstrb
	wire          hps_0_h2f_lw_axi_master_wready;                                 // mm_interconnect_1:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire   [11:0] hps_0_h2f_lw_axi_master_rid;                                    // mm_interconnect_1:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire          hps_0_h2f_lw_axi_master_rready;                                 // hps_0:h2f_lw_RREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_rready
	wire    [3:0] hps_0_h2f_lw_axi_master_awlen;                                  // hps_0:h2f_lw_AWLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlen
	wire   [11:0] hps_0_h2f_lw_axi_master_wid;                                    // hps_0:h2f_lw_WID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wid
	wire    [3:0] hps_0_h2f_lw_axi_master_arcache;                                // hps_0:h2f_lw_ARCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arcache
	wire          hps_0_h2f_lw_axi_master_wvalid;                                 // hps_0:h2f_lw_WVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wvalid
	wire   [20:0] hps_0_h2f_lw_axi_master_araddr;                                 // hps_0:h2f_lw_ARADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_araddr
	wire    [2:0] hps_0_h2f_lw_axi_master_arprot;                                 // hps_0:h2f_lw_ARPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arprot
	wire    [2:0] hps_0_h2f_lw_axi_master_awprot;                                 // hps_0:h2f_lw_AWPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awprot
	wire   [31:0] hps_0_h2f_lw_axi_master_wdata;                                  // hps_0:h2f_lw_WDATA -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wdata
	wire          hps_0_h2f_lw_axi_master_arvalid;                                // hps_0:h2f_lw_ARVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arvalid
	wire    [3:0] hps_0_h2f_lw_axi_master_awcache;                                // hps_0:h2f_lw_AWCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awcache
	wire   [11:0] hps_0_h2f_lw_axi_master_arid;                                   // hps_0:h2f_lw_ARID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arid
	wire    [1:0] hps_0_h2f_lw_axi_master_arlock;                                 // hps_0:h2f_lw_ARLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlock
	wire    [1:0] hps_0_h2f_lw_axi_master_awlock;                                 // hps_0:h2f_lw_AWLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlock
	wire   [20:0] hps_0_h2f_lw_axi_master_awaddr;                                 // hps_0:h2f_lw_AWADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awaddr
	wire    [1:0] hps_0_h2f_lw_axi_master_bresp;                                  // mm_interconnect_1:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire          hps_0_h2f_lw_axi_master_arready;                                // mm_interconnect_1:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire   [31:0] hps_0_h2f_lw_axi_master_rdata;                                  // mm_interconnect_1:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire          hps_0_h2f_lw_axi_master_awready;                                // mm_interconnect_1:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire    [1:0] hps_0_h2f_lw_axi_master_arburst;                                // hps_0:h2f_lw_ARBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arburst
	wire    [2:0] hps_0_h2f_lw_axi_master_arsize;                                 // hps_0:h2f_lw_ARSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arsize
	wire          hps_0_h2f_lw_axi_master_bready;                                 // hps_0:h2f_lw_BREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_bready
	wire          hps_0_h2f_lw_axi_master_rlast;                                  // mm_interconnect_1:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire          hps_0_h2f_lw_axi_master_wlast;                                  // hps_0:h2f_lw_WLAST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wlast
	wire    [1:0] hps_0_h2f_lw_axi_master_rresp;                                  // mm_interconnect_1:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire   [11:0] hps_0_h2f_lw_axi_master_awid;                                   // hps_0:h2f_lw_AWID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awid
	wire   [11:0] hps_0_h2f_lw_axi_master_bid;                                    // mm_interconnect_1:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire          hps_0_h2f_lw_axi_master_bvalid;                                 // mm_interconnect_1:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire    [2:0] hps_0_h2f_lw_axi_master_awsize;                                 // hps_0:h2f_lw_AWSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awsize
	wire          hps_0_h2f_lw_axi_master_awvalid;                                // hps_0:h2f_lw_AWVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awvalid
	wire          hps_0_h2f_lw_axi_master_rvalid;                                 // mm_interconnect_1:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire   [31:0] mm_interconnect_1_mm_bridge_lw_axi_s0_readdata;                 // mm_bridge_lw_axi:s0_readdata -> mm_interconnect_1:mm_bridge_lw_axi_s0_readdata
	wire          mm_interconnect_1_mm_bridge_lw_axi_s0_waitrequest;              // mm_bridge_lw_axi:s0_waitrequest -> mm_interconnect_1:mm_bridge_lw_axi_s0_waitrequest
	wire          mm_interconnect_1_mm_bridge_lw_axi_s0_debugaccess;              // mm_interconnect_1:mm_bridge_lw_axi_s0_debugaccess -> mm_bridge_lw_axi:s0_debugaccess
	wire   [14:0] mm_interconnect_1_mm_bridge_lw_axi_s0_address;                  // mm_interconnect_1:mm_bridge_lw_axi_s0_address -> mm_bridge_lw_axi:s0_address
	wire          mm_interconnect_1_mm_bridge_lw_axi_s0_read;                     // mm_interconnect_1:mm_bridge_lw_axi_s0_read -> mm_bridge_lw_axi:s0_read
	wire    [3:0] mm_interconnect_1_mm_bridge_lw_axi_s0_byteenable;               // mm_interconnect_1:mm_bridge_lw_axi_s0_byteenable -> mm_bridge_lw_axi:s0_byteenable
	wire          mm_interconnect_1_mm_bridge_lw_axi_s0_readdatavalid;            // mm_bridge_lw_axi:s0_readdatavalid -> mm_interconnect_1:mm_bridge_lw_axi_s0_readdatavalid
	wire          mm_interconnect_1_mm_bridge_lw_axi_s0_write;                    // mm_interconnect_1:mm_bridge_lw_axi_s0_write -> mm_bridge_lw_axi:s0_write
	wire   [31:0] mm_interconnect_1_mm_bridge_lw_axi_s0_writedata;                // mm_interconnect_1:mm_bridge_lw_axi_s0_writedata -> mm_bridge_lw_axi:s0_writedata
	wire    [0:0] mm_interconnect_1_mm_bridge_lw_axi_s0_burstcount;               // mm_interconnect_1:mm_bridge_lw_axi_s0_burstcount -> mm_bridge_lw_axi:s0_burstcount
	wire   [63:0] cnn_top_0_load_read_avalon_readdata;                            // mm_interconnect_2:cnn_top_0_load_read_avalon_readdata -> cnn_top_0:load_avm_readdata
	wire          cnn_top_0_load_read_avalon_waitrequest;                         // mm_interconnect_2:cnn_top_0_load_read_avalon_waitrequest -> cnn_top_0:load_avm_waitrequest
	wire   [31:0] cnn_top_0_load_read_avalon_address;                             // cnn_top_0:load_avm_address -> mm_interconnect_2:cnn_top_0_load_read_avalon_address
	wire    [7:0] cnn_top_0_load_read_avalon_byteenable;                          // cnn_top_0:load_avm_byteenable -> mm_interconnect_2:cnn_top_0_load_read_avalon_byteenable
	wire          cnn_top_0_load_read_avalon_read;                                // cnn_top_0:load_avm_read -> mm_interconnect_2:cnn_top_0_load_read_avalon_read
	wire          cnn_top_0_load_read_avalon_readdatavalid;                       // mm_interconnect_2:cnn_top_0_load_read_avalon_readdatavalid -> cnn_top_0:load_avm_readdatavalid
	wire    [4:0] cnn_top_0_load_read_avalon_burstcount;                          // cnn_top_0:load_avm_burstcount -> mm_interconnect_2:cnn_top_0_load_read_avalon_burstcount
	wire          cnn_top_0_output_read_avalon_waitrequest;                       // mm_interconnect_2:cnn_top_0_output_read_avalon_waitrequest -> cnn_top_0:output_avm_waitrequest
	wire   [31:0] cnn_top_0_output_read_avalon_address;                           // cnn_top_0:output_avm_address -> mm_interconnect_2:cnn_top_0_output_read_avalon_address
	wire    [7:0] cnn_top_0_output_read_avalon_byteenable;                        // cnn_top_0:output_avm_byteenable -> mm_interconnect_2:cnn_top_0_output_read_avalon_byteenable
	wire          cnn_top_0_output_read_avalon_write;                             // cnn_top_0:output_avm_write -> mm_interconnect_2:cnn_top_0_output_read_avalon_write
	wire   [63:0] cnn_top_0_output_read_avalon_writedata;                         // cnn_top_0:output_avm_writedata -> mm_interconnect_2:cnn_top_0_output_read_avalon_writedata
	wire    [4:0] cnn_top_0_output_read_avalon_burstcount;                        // cnn_top_0:output_avm_burstcount -> mm_interconnect_2:cnn_top_0_output_read_avalon_burstcount
	wire   [31:0] cnn_top_0_param_read_avalon_readdata;                           // mm_interconnect_2:cnn_top_0_param_read_avalon_readdata -> cnn_top_0:param_avm_readdata
	wire          cnn_top_0_param_read_avalon_waitrequest;                        // mm_interconnect_2:cnn_top_0_param_read_avalon_waitrequest -> cnn_top_0:param_avm_waitrequest
	wire   [31:0] cnn_top_0_param_read_avalon_address;                            // cnn_top_0:param_avm_address -> mm_interconnect_2:cnn_top_0_param_read_avalon_address
	wire    [3:0] cnn_top_0_param_read_avalon_byteenable;                         // cnn_top_0:param_avm_byteenable -> mm_interconnect_2:cnn_top_0_param_read_avalon_byteenable
	wire          cnn_top_0_param_read_avalon_read;                               // cnn_top_0:param_avm_read -> mm_interconnect_2:cnn_top_0_param_read_avalon_read
	wire          cnn_top_0_param_read_avalon_readdatavalid;                      // mm_interconnect_2:cnn_top_0_param_read_avalon_readdatavalid -> cnn_top_0:param_avm_readdatavalid
	wire    [4:0] cnn_top_0_param_read_avalon_burstcount;                         // cnn_top_0:param_avm_burstcount -> mm_interconnect_2:cnn_top_0_param_read_avalon_burstcount
	wire          cnn_top_0_scale_avm_avalon_waitrequest;                         // mm_interconnect_2:cnn_top_0_scale_avm_avalon_waitrequest -> cnn_top_0:scale_avm_waitrequest
	wire   [31:0] cnn_top_0_scale_avm_avalon_readdata;                            // mm_interconnect_2:cnn_top_0_scale_avm_avalon_readdata -> cnn_top_0:scale_avm_readdata
	wire   [31:0] cnn_top_0_scale_avm_avalon_address;                             // cnn_top_0:scale_avm_address -> mm_interconnect_2:cnn_top_0_scale_avm_avalon_address
	wire          cnn_top_0_scale_avm_avalon_read;                                // cnn_top_0:scale_avm_read -> mm_interconnect_2:cnn_top_0_scale_avm_avalon_read
	wire    [3:0] cnn_top_0_scale_avm_avalon_byteenable;                          // cnn_top_0:scale_avm_byteenable -> mm_interconnect_2:cnn_top_0_scale_avm_avalon_byteenable
	wire          cnn_top_0_scale_avm_avalon_readdatavalid;                       // mm_interconnect_2:cnn_top_0_scale_avm_avalon_readdatavalid -> cnn_top_0:scale_avm_readdatavalid
	wire    [4:0] cnn_top_0_scale_avm_avalon_burstcount;                          // cnn_top_0:scale_avm_burstcount -> mm_interconnect_2:cnn_top_0_scale_avm_avalon_burstcount
	wire  [127:0] mm_interconnect_2_mm_bridge_sdram0_s0_readdata;                 // mm_bridge_sdram0:s0_readdata -> mm_interconnect_2:mm_bridge_sdram0_s0_readdata
	wire          mm_interconnect_2_mm_bridge_sdram0_s0_waitrequest;              // mm_bridge_sdram0:s0_waitrequest -> mm_interconnect_2:mm_bridge_sdram0_s0_waitrequest
	wire          mm_interconnect_2_mm_bridge_sdram0_s0_debugaccess;              // mm_interconnect_2:mm_bridge_sdram0_s0_debugaccess -> mm_bridge_sdram0:s0_debugaccess
	wire   [31:0] mm_interconnect_2_mm_bridge_sdram0_s0_address;                  // mm_interconnect_2:mm_bridge_sdram0_s0_address -> mm_bridge_sdram0:s0_address
	wire          mm_interconnect_2_mm_bridge_sdram0_s0_read;                     // mm_interconnect_2:mm_bridge_sdram0_s0_read -> mm_bridge_sdram0:s0_read
	wire   [15:0] mm_interconnect_2_mm_bridge_sdram0_s0_byteenable;               // mm_interconnect_2:mm_bridge_sdram0_s0_byteenable -> mm_bridge_sdram0:s0_byteenable
	wire          mm_interconnect_2_mm_bridge_sdram0_s0_readdatavalid;            // mm_bridge_sdram0:s0_readdatavalid -> mm_interconnect_2:mm_bridge_sdram0_s0_readdatavalid
	wire          mm_interconnect_2_mm_bridge_sdram0_s0_write;                    // mm_interconnect_2:mm_bridge_sdram0_s0_write -> mm_bridge_sdram0:s0_write
	wire  [127:0] mm_interconnect_2_mm_bridge_sdram0_s0_writedata;                // mm_interconnect_2:mm_bridge_sdram0_s0_writedata -> mm_bridge_sdram0:s0_writedata
	wire    [4:0] mm_interconnect_2_mm_bridge_sdram0_s0_burstcount;               // mm_interconnect_2:mm_bridge_sdram0_s0_burstcount -> mm_bridge_sdram0:s0_burstcount
	wire          mm_bridge_lw_axi_m0_waitrequest;                                // mm_interconnect_3:mm_bridge_lw_axi_m0_waitrequest -> mm_bridge_lw_axi:m0_waitrequest
	wire   [31:0] mm_bridge_lw_axi_m0_readdata;                                   // mm_interconnect_3:mm_bridge_lw_axi_m0_readdata -> mm_bridge_lw_axi:m0_readdata
	wire          mm_bridge_lw_axi_m0_debugaccess;                                // mm_bridge_lw_axi:m0_debugaccess -> mm_interconnect_3:mm_bridge_lw_axi_m0_debugaccess
	wire   [14:0] mm_bridge_lw_axi_m0_address;                                    // mm_bridge_lw_axi:m0_address -> mm_interconnect_3:mm_bridge_lw_axi_m0_address
	wire          mm_bridge_lw_axi_m0_read;                                       // mm_bridge_lw_axi:m0_read -> mm_interconnect_3:mm_bridge_lw_axi_m0_read
	wire    [3:0] mm_bridge_lw_axi_m0_byteenable;                                 // mm_bridge_lw_axi:m0_byteenable -> mm_interconnect_3:mm_bridge_lw_axi_m0_byteenable
	wire          mm_bridge_lw_axi_m0_readdatavalid;                              // mm_interconnect_3:mm_bridge_lw_axi_m0_readdatavalid -> mm_bridge_lw_axi:m0_readdatavalid
	wire   [31:0] mm_bridge_lw_axi_m0_writedata;                                  // mm_bridge_lw_axi:m0_writedata -> mm_interconnect_3:mm_bridge_lw_axi_m0_writedata
	wire          mm_bridge_lw_axi_m0_write;                                      // mm_bridge_lw_axi:m0_write -> mm_interconnect_3:mm_bridge_lw_axi_m0_write
	wire    [0:0] mm_bridge_lw_axi_m0_burstcount;                                 // mm_bridge_lw_axi:m0_burstcount -> mm_interconnect_3:mm_bridge_lw_axi_m0_burstcount
	wire   [31:0] fpga_only_master_master_readdata;                               // mm_interconnect_3:fpga_only_master_master_readdata -> fpga_only_master:master_readdata
	wire          fpga_only_master_master_waitrequest;                            // mm_interconnect_3:fpga_only_master_master_waitrequest -> fpga_only_master:master_waitrequest
	wire   [31:0] fpga_only_master_master_address;                                // fpga_only_master:master_address -> mm_interconnect_3:fpga_only_master_master_address
	wire          fpga_only_master_master_read;                                   // fpga_only_master:master_read -> mm_interconnect_3:fpga_only_master_master_read
	wire    [3:0] fpga_only_master_master_byteenable;                             // fpga_only_master:master_byteenable -> mm_interconnect_3:fpga_only_master_master_byteenable
	wire          fpga_only_master_master_readdatavalid;                          // mm_interconnect_3:fpga_only_master_master_readdatavalid -> fpga_only_master:master_readdatavalid
	wire          fpga_only_master_master_write;                                  // fpga_only_master:master_write -> mm_interconnect_3:fpga_only_master_master_write
	wire   [31:0] fpga_only_master_master_writedata;                              // fpga_only_master:master_writedata -> mm_interconnect_3:fpga_only_master_master_writedata
	wire   [31:0] mm_interconnect_3_vcam_0_cfg_bus_readdata;                      // vcam_0:cfg_read_data -> mm_interconnect_3:vcam_0_cfg_bus_readdata
	wire    [3:0] mm_interconnect_3_vcam_0_cfg_bus_address;                       // mm_interconnect_3:vcam_0_cfg_bus_address -> vcam_0:cfg_addr
	wire          mm_interconnect_3_vcam_0_cfg_bus_read;                          // mm_interconnect_3:vcam_0_cfg_bus_read -> vcam_0:cfg_read
	wire          mm_interconnect_3_vcam_0_cfg_bus_write;                         // mm_interconnect_3:vcam_0_cfg_bus_write -> vcam_0:cfg_write
	wire   [31:0] mm_interconnect_3_vcam_0_cfg_bus_writedata;                     // mm_interconnect_3:vcam_0_cfg_bus_writedata -> vcam_0:cfg_write_data
	wire   [31:0] mm_interconnect_3_dvp_ddr3_0_cfg_bus_readdata;                  // dvp_ddr3_0:avalon_read_data -> mm_interconnect_3:dvp_ddr3_0_cfg_bus_readdata
	wire    [3:0] mm_interconnect_3_dvp_ddr3_0_cfg_bus_address;                   // mm_interconnect_3:dvp_ddr3_0_cfg_bus_address -> dvp_ddr3_0:avalon_addr
	wire          mm_interconnect_3_dvp_ddr3_0_cfg_bus_read;                      // mm_interconnect_3:dvp_ddr3_0_cfg_bus_read -> dvp_ddr3_0:avalon_read
	wire          mm_interconnect_3_dvp_ddr3_0_cfg_bus_write;                     // mm_interconnect_3:dvp_ddr3_0_cfg_bus_write -> dvp_ddr3_0:avalon_write
	wire   [31:0] mm_interconnect_3_dvp_ddr3_0_cfg_bus_writedata;                 // mm_interconnect_3:dvp_ddr3_0_cfg_bus_writedata -> dvp_ddr3_0:avalon_write_data
	wire   [31:0] mm_interconnect_3_ddr3_vga_0_cfg_bus_readdata;                  // ddr3_vga_0:avalon_read_data -> mm_interconnect_3:ddr3_vga_0_cfg_bus_readdata
	wire    [3:0] mm_interconnect_3_ddr3_vga_0_cfg_bus_address;                   // mm_interconnect_3:ddr3_vga_0_cfg_bus_address -> ddr3_vga_0:avalon_addr
	wire          mm_interconnect_3_ddr3_vga_0_cfg_bus_read;                      // mm_interconnect_3:ddr3_vga_0_cfg_bus_read -> ddr3_vga_0:avalon_read
	wire          mm_interconnect_3_ddr3_vga_0_cfg_bus_write;                     // mm_interconnect_3:ddr3_vga_0_cfg_bus_write -> ddr3_vga_0:avalon_write
	wire   [31:0] mm_interconnect_3_ddr3_vga_0_cfg_bus_writedata;                 // mm_interconnect_3:ddr3_vga_0_cfg_bus_writedata -> ddr3_vga_0:avalon_write_data
	wire   [31:0] mm_interconnect_3_sysid_qsys_control_slave_readdata;            // sysid_qsys:readdata -> mm_interconnect_3:sysid_qsys_control_slave_readdata
	wire    [0:0] mm_interconnect_3_sysid_qsys_control_slave_address;             // mm_interconnect_3:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire   [31:0] mm_interconnect_3_cnn_top_0_hps2cnn_avs_readdata;               // cnn_top_0:as_readdata -> mm_interconnect_3:cnn_top_0_hps2cnn_avs_readdata
	wire          mm_interconnect_3_cnn_top_0_hps2cnn_avs_waitrequest;            // cnn_top_0:as_data_waitquest -> mm_interconnect_3:cnn_top_0_hps2cnn_avs_waitrequest
	wire    [7:0] mm_interconnect_3_cnn_top_0_hps2cnn_avs_address;                // mm_interconnect_3:cnn_top_0_hps2cnn_avs_address -> cnn_top_0:as_address
	wire          mm_interconnect_3_cnn_top_0_hps2cnn_avs_read;                   // mm_interconnect_3:cnn_top_0_hps2cnn_avs_read -> cnn_top_0:as_read
	wire          mm_interconnect_3_cnn_top_0_hps2cnn_avs_write;                  // mm_interconnect_3:cnn_top_0_hps2cnn_avs_write -> cnn_top_0:as_write
	wire   [31:0] mm_interconnect_3_cnn_top_0_hps2cnn_avs_writedata;              // mm_interconnect_3:cnn_top_0_hps2cnn_avs_writedata -> cnn_top_0:as_writedata
	wire   [31:0] mm_interconnect_3_sld_hub_controller_system_0_s0_readdata;      // sld_hub_controller_system_0:s0_readdata -> mm_interconnect_3:sld_hub_controller_system_0_s0_readdata
	wire          mm_interconnect_3_sld_hub_controller_system_0_s0_waitrequest;   // sld_hub_controller_system_0:s0_waitrequest -> mm_interconnect_3:sld_hub_controller_system_0_s0_waitrequest
	wire          mm_interconnect_3_sld_hub_controller_system_0_s0_debugaccess;   // mm_interconnect_3:sld_hub_controller_system_0_s0_debugaccess -> sld_hub_controller_system_0:s0_debugaccess
	wire    [6:0] mm_interconnect_3_sld_hub_controller_system_0_s0_address;       // mm_interconnect_3:sld_hub_controller_system_0_s0_address -> sld_hub_controller_system_0:s0_address
	wire          mm_interconnect_3_sld_hub_controller_system_0_s0_read;          // mm_interconnect_3:sld_hub_controller_system_0_s0_read -> sld_hub_controller_system_0:s0_read
	wire    [3:0] mm_interconnect_3_sld_hub_controller_system_0_s0_byteenable;    // mm_interconnect_3:sld_hub_controller_system_0_s0_byteenable -> sld_hub_controller_system_0:s0_byteenable
	wire          mm_interconnect_3_sld_hub_controller_system_0_s0_readdatavalid; // sld_hub_controller_system_0:s0_readdatavalid -> mm_interconnect_3:sld_hub_controller_system_0_s0_readdatavalid
	wire          mm_interconnect_3_sld_hub_controller_system_0_s0_write;         // mm_interconnect_3:sld_hub_controller_system_0_s0_write -> sld_hub_controller_system_0:s0_write
	wire   [31:0] mm_interconnect_3_sld_hub_controller_system_0_s0_writedata;     // mm_interconnect_3:sld_hub_controller_system_0_s0_writedata -> sld_hub_controller_system_0:s0_writedata
	wire    [0:0] mm_interconnect_3_sld_hub_controller_system_0_s0_burstcount;    // mm_interconnect_3:sld_hub_controller_system_0_s0_burstcount -> sld_hub_controller_system_0:s0_burstcount
	wire          mm_interconnect_3_button_pio_s1_chipselect;                     // mm_interconnect_3:button_pio_s1_chipselect -> button_pio:chipselect
	wire   [31:0] mm_interconnect_3_button_pio_s1_readdata;                       // button_pio:readdata -> mm_interconnect_3:button_pio_s1_readdata
	wire    [1:0] mm_interconnect_3_button_pio_s1_address;                        // mm_interconnect_3:button_pio_s1_address -> button_pio:address
	wire          mm_interconnect_3_button_pio_s1_write;                          // mm_interconnect_3:button_pio_s1_write -> button_pio:write_n
	wire   [31:0] mm_interconnect_3_button_pio_s1_writedata;                      // mm_interconnect_3:button_pio_s1_writedata -> button_pio:writedata
	wire          mm_interconnect_3_dipsw_pio_s1_chipselect;                      // mm_interconnect_3:dipsw_pio_s1_chipselect -> dipsw_pio:chipselect
	wire   [31:0] mm_interconnect_3_dipsw_pio_s1_readdata;                        // dipsw_pio:readdata -> mm_interconnect_3:dipsw_pio_s1_readdata
	wire    [1:0] mm_interconnect_3_dipsw_pio_s1_address;                         // mm_interconnect_3:dipsw_pio_s1_address -> dipsw_pio:address
	wire          mm_interconnect_3_dipsw_pio_s1_write;                           // mm_interconnect_3:dipsw_pio_s1_write -> dipsw_pio:write_n
	wire   [31:0] mm_interconnect_3_dipsw_pio_s1_writedata;                       // mm_interconnect_3:dipsw_pio_s1_writedata -> dipsw_pio:writedata
	wire          mm_interconnect_3_led_pio_s1_chipselect;                        // mm_interconnect_3:led_pio_s1_chipselect -> led_pio:chipselect
	wire   [31:0] mm_interconnect_3_led_pio_s1_readdata;                          // led_pio:readdata -> mm_interconnect_3:led_pio_s1_readdata
	wire    [1:0] mm_interconnect_3_led_pio_s1_address;                           // mm_interconnect_3:led_pio_s1_address -> led_pio:address
	wire          mm_interconnect_3_led_pio_s1_write;                             // mm_interconnect_3:led_pio_s1_write -> led_pio:write_n
	wire   [31:0] mm_interconnect_3_led_pio_s1_writedata;                         // mm_interconnect_3:led_pio_s1_writedata -> led_pio:writedata
	wire          mm_interconnect_3_vhdmi_0_s_avalon_mm_chipselect;               // mm_interconnect_3:vhdmi_0_s_avalon_mm_chipselect -> vhdmi_0:s_avl_chipselect
	wire   [31:0] mm_interconnect_3_vhdmi_0_s_avalon_mm_readdata;                 // vhdmi_0:s_avl_rd_data -> mm_interconnect_3:vhdmi_0_s_avalon_mm_readdata
	wire    [7:0] mm_interconnect_3_vhdmi_0_s_avalon_mm_address;                  // mm_interconnect_3:vhdmi_0_s_avalon_mm_address -> vhdmi_0:s_avl_address
	wire          mm_interconnect_3_vhdmi_0_s_avalon_mm_read;                     // mm_interconnect_3:vhdmi_0_s_avalon_mm_read -> vhdmi_0:s_avl_rd_req
	wire          mm_interconnect_3_vhdmi_0_s_avalon_mm_write;                    // mm_interconnect_3:vhdmi_0_s_avalon_mm_write -> vhdmi_0:s_avl_wr_req
	wire   [31:0] mm_interconnect_3_vhdmi_0_s_avalon_mm_writedata;                // mm_interconnect_3:vhdmi_0_s_avalon_mm_writedata -> vhdmi_0:s_avl_wr_data
	wire          mm_bridge_axi_m0_waitrequest;                                   // mm_interconnect_4:mm_bridge_axi_m0_waitrequest -> mm_bridge_axi:m0_waitrequest
	wire  [127:0] mm_bridge_axi_m0_readdata;                                      // mm_interconnect_4:mm_bridge_axi_m0_readdata -> mm_bridge_axi:m0_readdata
	wire          mm_bridge_axi_m0_debugaccess;                                   // mm_bridge_axi:m0_debugaccess -> mm_interconnect_4:mm_bridge_axi_m0_debugaccess
	wire   [31:0] mm_bridge_axi_m0_address;                                       // mm_bridge_axi:m0_address -> mm_interconnect_4:mm_bridge_axi_m0_address
	wire          mm_bridge_axi_m0_read;                                          // mm_bridge_axi:m0_read -> mm_interconnect_4:mm_bridge_axi_m0_read
	wire   [15:0] mm_bridge_axi_m0_byteenable;                                    // mm_bridge_axi:m0_byteenable -> mm_interconnect_4:mm_bridge_axi_m0_byteenable
	wire          mm_bridge_axi_m0_readdatavalid;                                 // mm_interconnect_4:mm_bridge_axi_m0_readdatavalid -> mm_bridge_axi:m0_readdatavalid
	wire  [127:0] mm_bridge_axi_m0_writedata;                                     // mm_bridge_axi:m0_writedata -> mm_interconnect_4:mm_bridge_axi_m0_writedata
	wire          mm_bridge_axi_m0_write;                                         // mm_bridge_axi:m0_write -> mm_interconnect_4:mm_bridge_axi_m0_write
	wire    [4:0] mm_bridge_axi_m0_burstcount;                                    // mm_bridge_axi:m0_burstcount -> mm_interconnect_4:mm_bridge_axi_m0_burstcount
	wire   [31:0] hps_only_master_master_readdata;                                // mm_interconnect_4:hps_only_master_master_readdata -> hps_only_master:master_readdata
	wire          hps_only_master_master_waitrequest;                             // mm_interconnect_4:hps_only_master_master_waitrequest -> hps_only_master:master_waitrequest
	wire   [31:0] hps_only_master_master_address;                                 // hps_only_master:master_address -> mm_interconnect_4:hps_only_master_master_address
	wire          hps_only_master_master_read;                                    // hps_only_master:master_read -> mm_interconnect_4:hps_only_master_master_read
	wire    [3:0] hps_only_master_master_byteenable;                              // hps_only_master:master_byteenable -> mm_interconnect_4:hps_only_master_master_byteenable
	wire          hps_only_master_master_readdatavalid;                           // mm_interconnect_4:hps_only_master_master_readdatavalid -> hps_only_master:master_readdatavalid
	wire          hps_only_master_master_write;                                   // hps_only_master:master_write -> mm_interconnect_4:hps_only_master_master_write
	wire   [31:0] hps_only_master_master_writedata;                               // hps_only_master:master_writedata -> mm_interconnect_4:hps_only_master_master_writedata
	wire    [1:0] mm_interconnect_4_hps_0_f2h_axi_slave_awburst;                  // mm_interconnect_4:hps_0_f2h_axi_slave_awburst -> hps_0:f2h_AWBURST
	wire    [4:0] mm_interconnect_4_hps_0_f2h_axi_slave_awuser;                   // mm_interconnect_4:hps_0_f2h_axi_slave_awuser -> hps_0:f2h_AWUSER
	wire    [3:0] mm_interconnect_4_hps_0_f2h_axi_slave_arlen;                    // mm_interconnect_4:hps_0_f2h_axi_slave_arlen -> hps_0:f2h_ARLEN
	wire   [15:0] mm_interconnect_4_hps_0_f2h_axi_slave_wstrb;                    // mm_interconnect_4:hps_0_f2h_axi_slave_wstrb -> hps_0:f2h_WSTRB
	wire          mm_interconnect_4_hps_0_f2h_axi_slave_wready;                   // hps_0:f2h_WREADY -> mm_interconnect_4:hps_0_f2h_axi_slave_wready
	wire    [7:0] mm_interconnect_4_hps_0_f2h_axi_slave_rid;                      // hps_0:f2h_RID -> mm_interconnect_4:hps_0_f2h_axi_slave_rid
	wire          mm_interconnect_4_hps_0_f2h_axi_slave_rready;                   // mm_interconnect_4:hps_0_f2h_axi_slave_rready -> hps_0:f2h_RREADY
	wire    [3:0] mm_interconnect_4_hps_0_f2h_axi_slave_awlen;                    // mm_interconnect_4:hps_0_f2h_axi_slave_awlen -> hps_0:f2h_AWLEN
	wire    [7:0] mm_interconnect_4_hps_0_f2h_axi_slave_wid;                      // mm_interconnect_4:hps_0_f2h_axi_slave_wid -> hps_0:f2h_WID
	wire    [3:0] mm_interconnect_4_hps_0_f2h_axi_slave_arcache;                  // mm_interconnect_4:hps_0_f2h_axi_slave_arcache -> hps_0:f2h_ARCACHE
	wire          mm_interconnect_4_hps_0_f2h_axi_slave_wvalid;                   // mm_interconnect_4:hps_0_f2h_axi_slave_wvalid -> hps_0:f2h_WVALID
	wire   [31:0] mm_interconnect_4_hps_0_f2h_axi_slave_araddr;                   // mm_interconnect_4:hps_0_f2h_axi_slave_araddr -> hps_0:f2h_ARADDR
	wire    [2:0] mm_interconnect_4_hps_0_f2h_axi_slave_arprot;                   // mm_interconnect_4:hps_0_f2h_axi_slave_arprot -> hps_0:f2h_ARPROT
	wire    [2:0] mm_interconnect_4_hps_0_f2h_axi_slave_awprot;                   // mm_interconnect_4:hps_0_f2h_axi_slave_awprot -> hps_0:f2h_AWPROT
	wire  [127:0] mm_interconnect_4_hps_0_f2h_axi_slave_wdata;                    // mm_interconnect_4:hps_0_f2h_axi_slave_wdata -> hps_0:f2h_WDATA
	wire          mm_interconnect_4_hps_0_f2h_axi_slave_arvalid;                  // mm_interconnect_4:hps_0_f2h_axi_slave_arvalid -> hps_0:f2h_ARVALID
	wire    [3:0] mm_interconnect_4_hps_0_f2h_axi_slave_awcache;                  // mm_interconnect_4:hps_0_f2h_axi_slave_awcache -> hps_0:f2h_AWCACHE
	wire    [7:0] mm_interconnect_4_hps_0_f2h_axi_slave_arid;                     // mm_interconnect_4:hps_0_f2h_axi_slave_arid -> hps_0:f2h_ARID
	wire    [1:0] mm_interconnect_4_hps_0_f2h_axi_slave_arlock;                   // mm_interconnect_4:hps_0_f2h_axi_slave_arlock -> hps_0:f2h_ARLOCK
	wire    [1:0] mm_interconnect_4_hps_0_f2h_axi_slave_awlock;                   // mm_interconnect_4:hps_0_f2h_axi_slave_awlock -> hps_0:f2h_AWLOCK
	wire   [31:0] mm_interconnect_4_hps_0_f2h_axi_slave_awaddr;                   // mm_interconnect_4:hps_0_f2h_axi_slave_awaddr -> hps_0:f2h_AWADDR
	wire    [1:0] mm_interconnect_4_hps_0_f2h_axi_slave_bresp;                    // hps_0:f2h_BRESP -> mm_interconnect_4:hps_0_f2h_axi_slave_bresp
	wire          mm_interconnect_4_hps_0_f2h_axi_slave_arready;                  // hps_0:f2h_ARREADY -> mm_interconnect_4:hps_0_f2h_axi_slave_arready
	wire  [127:0] mm_interconnect_4_hps_0_f2h_axi_slave_rdata;                    // hps_0:f2h_RDATA -> mm_interconnect_4:hps_0_f2h_axi_slave_rdata
	wire          mm_interconnect_4_hps_0_f2h_axi_slave_awready;                  // hps_0:f2h_AWREADY -> mm_interconnect_4:hps_0_f2h_axi_slave_awready
	wire    [1:0] mm_interconnect_4_hps_0_f2h_axi_slave_arburst;                  // mm_interconnect_4:hps_0_f2h_axi_slave_arburst -> hps_0:f2h_ARBURST
	wire    [2:0] mm_interconnect_4_hps_0_f2h_axi_slave_arsize;                   // mm_interconnect_4:hps_0_f2h_axi_slave_arsize -> hps_0:f2h_ARSIZE
	wire          mm_interconnect_4_hps_0_f2h_axi_slave_bready;                   // mm_interconnect_4:hps_0_f2h_axi_slave_bready -> hps_0:f2h_BREADY
	wire          mm_interconnect_4_hps_0_f2h_axi_slave_rlast;                    // hps_0:f2h_RLAST -> mm_interconnect_4:hps_0_f2h_axi_slave_rlast
	wire          mm_interconnect_4_hps_0_f2h_axi_slave_wlast;                    // mm_interconnect_4:hps_0_f2h_axi_slave_wlast -> hps_0:f2h_WLAST
	wire    [1:0] mm_interconnect_4_hps_0_f2h_axi_slave_rresp;                    // hps_0:f2h_RRESP -> mm_interconnect_4:hps_0_f2h_axi_slave_rresp
	wire    [7:0] mm_interconnect_4_hps_0_f2h_axi_slave_awid;                     // mm_interconnect_4:hps_0_f2h_axi_slave_awid -> hps_0:f2h_AWID
	wire    [7:0] mm_interconnect_4_hps_0_f2h_axi_slave_bid;                      // hps_0:f2h_BID -> mm_interconnect_4:hps_0_f2h_axi_slave_bid
	wire          mm_interconnect_4_hps_0_f2h_axi_slave_bvalid;                   // hps_0:f2h_BVALID -> mm_interconnect_4:hps_0_f2h_axi_slave_bvalid
	wire    [2:0] mm_interconnect_4_hps_0_f2h_axi_slave_awsize;                   // mm_interconnect_4:hps_0_f2h_axi_slave_awsize -> hps_0:f2h_AWSIZE
	wire          mm_interconnect_4_hps_0_f2h_axi_slave_awvalid;                  // mm_interconnect_4:hps_0_f2h_axi_slave_awvalid -> hps_0:f2h_AWVALID
	wire    [4:0] mm_interconnect_4_hps_0_f2h_axi_slave_aruser;                   // mm_interconnect_4:hps_0_f2h_axi_slave_aruser -> hps_0:f2h_ARUSER
	wire          mm_interconnect_4_hps_0_f2h_axi_slave_rvalid;                   // hps_0:f2h_RVALID -> mm_interconnect_4:hps_0_f2h_axi_slave_rvalid
	wire          mm_bridge_sdram0_m0_waitrequest;                                // mm_interconnect_5:mm_bridge_sdram0_m0_waitrequest -> mm_bridge_sdram0:m0_waitrequest
	wire  [127:0] mm_bridge_sdram0_m0_readdata;                                   // mm_interconnect_5:mm_bridge_sdram0_m0_readdata -> mm_bridge_sdram0:m0_readdata
	wire          mm_bridge_sdram0_m0_debugaccess;                                // mm_bridge_sdram0:m0_debugaccess -> mm_interconnect_5:mm_bridge_sdram0_m0_debugaccess
	wire   [31:0] mm_bridge_sdram0_m0_address;                                    // mm_bridge_sdram0:m0_address -> mm_interconnect_5:mm_bridge_sdram0_m0_address
	wire          mm_bridge_sdram0_m0_read;                                       // mm_bridge_sdram0:m0_read -> mm_interconnect_5:mm_bridge_sdram0_m0_read
	wire   [15:0] mm_bridge_sdram0_m0_byteenable;                                 // mm_bridge_sdram0:m0_byteenable -> mm_interconnect_5:mm_bridge_sdram0_m0_byteenable
	wire          mm_bridge_sdram0_m0_readdatavalid;                              // mm_interconnect_5:mm_bridge_sdram0_m0_readdatavalid -> mm_bridge_sdram0:m0_readdatavalid
	wire  [127:0] mm_bridge_sdram0_m0_writedata;                                  // mm_bridge_sdram0:m0_writedata -> mm_interconnect_5:mm_bridge_sdram0_m0_writedata
	wire          mm_bridge_sdram0_m0_write;                                      // mm_bridge_sdram0:m0_write -> mm_interconnect_5:mm_bridge_sdram0_m0_write
	wire    [4:0] mm_bridge_sdram0_m0_burstcount;                                 // mm_bridge_sdram0:m0_burstcount -> mm_interconnect_5:mm_bridge_sdram0_m0_burstcount
	wire   [31:0] f2sdram_only_master_master_readdata;                            // mm_interconnect_5:f2sdram_only_master_master_readdata -> f2sdram_only_master:master_readdata
	wire          f2sdram_only_master_master_waitrequest;                         // mm_interconnect_5:f2sdram_only_master_master_waitrequest -> f2sdram_only_master:master_waitrequest
	wire   [31:0] f2sdram_only_master_master_address;                             // f2sdram_only_master:master_address -> mm_interconnect_5:f2sdram_only_master_master_address
	wire          f2sdram_only_master_master_read;                                // f2sdram_only_master:master_read -> mm_interconnect_5:f2sdram_only_master_master_read
	wire    [3:0] f2sdram_only_master_master_byteenable;                          // f2sdram_only_master:master_byteenable -> mm_interconnect_5:f2sdram_only_master_master_byteenable
	wire          f2sdram_only_master_master_readdatavalid;                       // mm_interconnect_5:f2sdram_only_master_master_readdatavalid -> f2sdram_only_master:master_readdatavalid
	wire          f2sdram_only_master_master_write;                               // f2sdram_only_master:master_write -> mm_interconnect_5:f2sdram_only_master_master_write
	wire   [31:0] f2sdram_only_master_master_writedata;                           // f2sdram_only_master:master_writedata -> mm_interconnect_5:f2sdram_only_master_master_writedata
	wire  [127:0] mm_interconnect_5_hps_0_f2h_sdram0_data_readdata;               // hps_0:f2h_sdram0_READDATA -> mm_interconnect_5:hps_0_f2h_sdram0_data_readdata
	wire          mm_interconnect_5_hps_0_f2h_sdram0_data_waitrequest;            // hps_0:f2h_sdram0_WAITREQUEST -> mm_interconnect_5:hps_0_f2h_sdram0_data_waitrequest
	wire   [27:0] mm_interconnect_5_hps_0_f2h_sdram0_data_address;                // mm_interconnect_5:hps_0_f2h_sdram0_data_address -> hps_0:f2h_sdram0_ADDRESS
	wire          mm_interconnect_5_hps_0_f2h_sdram0_data_read;                   // mm_interconnect_5:hps_0_f2h_sdram0_data_read -> hps_0:f2h_sdram0_READ
	wire   [15:0] mm_interconnect_5_hps_0_f2h_sdram0_data_byteenable;             // mm_interconnect_5:hps_0_f2h_sdram0_data_byteenable -> hps_0:f2h_sdram0_BYTEENABLE
	wire          mm_interconnect_5_hps_0_f2h_sdram0_data_readdatavalid;          // hps_0:f2h_sdram0_READDATAVALID -> mm_interconnect_5:hps_0_f2h_sdram0_data_readdatavalid
	wire          mm_interconnect_5_hps_0_f2h_sdram0_data_write;                  // mm_interconnect_5:hps_0_f2h_sdram0_data_write -> hps_0:f2h_sdram0_WRITE
	wire  [127:0] mm_interconnect_5_hps_0_f2h_sdram0_data_writedata;              // mm_interconnect_5:hps_0_f2h_sdram0_data_writedata -> hps_0:f2h_sdram0_WRITEDATA
	wire    [7:0] mm_interconnect_5_hps_0_f2h_sdram0_data_burstcount;             // mm_interconnect_5:hps_0_f2h_sdram0_data_burstcount -> hps_0:f2h_sdram0_BURSTCOUNT
	wire   [31:0] hps_0_f2h_irq0_irq;                                             // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire   [31:0] hps_0_f2h_irq1_irq;                                             // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire          rst_controller_reset_out_reset;                                 // rst_controller:reset_out -> [button_pio:reset_n, ddr3_vga_0:rst_n, dipsw_pio:reset_n, dvp_ddr3_0:rst_n, led_pio:reset_n, mm_bridge_axi:reset, mm_bridge_lw_axi:reset, mm_interconnect_0:vcam_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:mm_bridge_lw_axi_reset_reset_bridge_in_reset_reset, mm_interconnect_3:fpga_only_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_3:mm_bridge_lw_axi_reset_reset_bridge_in_reset_reset, mm_interconnect_4:hps_only_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_4:mm_bridge_axi_reset_reset_bridge_in_reset_reset, mm_interconnect_5:f2sdram_only_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_5:f2sdram_only_master_master_translator_reset_reset_bridge_in_reset_reset, sld_hub_controller_system_0:reset_reset, sysid_qsys:reset_n, vcam_0:rst_n, vhdmi_0:rst_n]
	wire          rst_controller_001_reset_out_reset;                             // rst_controller_001:reset_out -> [cnn_top_0:rst_n, mm_bridge_sdram0:reset, mm_interconnect_2:cnn_top_0_reset_reset_bridge_in_reset_reset, mm_interconnect_3:cnn_top_0_reset_reset_bridge_in_reset_reset, mm_interconnect_5:mm_bridge_sdram0_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_002_reset_out_reset;                             // rst_controller_002:reset_out -> [mm_interconnect_1:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_4:hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset]
	wire          rst_controller_003_reset_out_reset;                             // rst_controller_003:reset_out -> mm_interconnect_5:hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset

	soc_system_button_pio button_pio (
		.clk        (clk_50_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_3_button_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_3_button_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_3_button_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_3_button_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_3_button_pio_s1_readdata),   //                    .readdata
		.out_port   (button_pio_external_connection_export)       // external_connection.export
	);

	cnn_top #(
		.OUTPUT_CHANNEL_TILE     (8),
		.INPUT_CHANNEL_TILE      (8),
		.INPUT_WIDTH             (8),
		.WEIGHT_WIDTH            (8),
		.INPUT_ROW_TILE          (11),
		.IMAGE_MAX_W             (302),
		.OUTPUT_ROW_TILE         (5),
		.OUTPUT_MAX_W            (150),
		.IN_C_WIDTH              (11),
		.IN_H_WIDTH              (9),
		.IN_W_WIDTH              (9),
		.OUTPUT_C_WIDTH          (11),
		.OUTPUT_H_WIDTH          (9),
		.OUTPUT_W_WIDTH          (9),
		.KERNEL_WIDTH            (2),
		.KERNEL_SIZE_WIDTH       (4),
		.INPUT_PAD_WIDTH         (2),
		.OUTPUT_PAD_WIDTH        (2),
		.CNN_TYPE_WIDTH          (3),
		.CNN_STRIDE_WIDTH        (2),
		.CNN_RELU_WIDTH          (3),
		.KERNAL_SIZE             (9),
		.CFG_PARAM_WIDTH         (32),
		.OUTPUT_ADDR_WIDTH       (10),
		.OUTPUT_WIDTH            (32),
		.SCALE_6                 (34'b0001000000110000000000000000000000),
		.REORGANIZE_BUFF_DEEP    (2048),
		.REORG_RAM_ADDR_WIDTH    (7),
		.REORG_RAM_DATA_WIDTH    (128),
		.REORG_RAM_SEL_WIDTH     (16),
		.INPUT_RAM_DATA_WIDTH    (64),
		.CFG_M_AXI_ADDR_WIDTH    (32),
		.CFG_M_AXI_DATA_WIDTH    (32),
		.LOAD_M_AXI_ADDR_WIDTH   (32),
		.LOAD_M_AXI_DATA_WIDTH   (64),
		.REORG_M_AXI_ADDR_WIDTH  (32),
		.REORG_M_AXI_DATA_WIDTH  (8),
		.SCALE_M_AXI_ADDR_WIDTH  (32),
		.SCALE_M_AXI_DATA_WIDTH  (32),
		.OUTPUT_M_AXI_ADDR_WIDTH (32),
		.OUTPUT_M_AXI_DATA_WIDTH (64)
	) cnn_top_0 (
		.rst_n                   (~rst_controller_001_reset_out_reset),                 //              reset.reset_n
		.as_address              (mm_interconnect_3_cnn_top_0_hps2cnn_avs_address),     //        hps2cnn_avs.address
		.as_write                (mm_interconnect_3_cnn_top_0_hps2cnn_avs_write),       //                   .write
		.as_read                 (mm_interconnect_3_cnn_top_0_hps2cnn_avs_read),        //                   .read
		.as_writedata            (mm_interconnect_3_cnn_top_0_hps2cnn_avs_writedata),   //                   .writedata
		.as_readdata             (mm_interconnect_3_cnn_top_0_hps2cnn_avs_readdata),    //                   .readdata
		.as_data_waitquest       (mm_interconnect_3_cnn_top_0_hps2cnn_avs_waitrequest), //                   .waitrequest
		.sysclk                  (clk_cnn_clk),                                         //            clock_1.clk
		.param_avm_address       (cnn_top_0_param_read_avalon_address),                 //  param_read_avalon.address
		.param_avm_burstcount    (cnn_top_0_param_read_avalon_burstcount),              //                   .burstcount
		.param_avm_byteenable    (cnn_top_0_param_read_avalon_byteenable),              //                   .byteenable
		.param_avm_read          (cnn_top_0_param_read_avalon_read),                    //                   .read
		.param_avm_readdata      (cnn_top_0_param_read_avalon_readdata),                //                   .readdata
		.param_avm_readdatavalid (cnn_top_0_param_read_avalon_readdatavalid),           //                   .readdatavalid
		.param_avm_waitrequest   (cnn_top_0_param_read_avalon_waitrequest),             //                   .waitrequest
		.load_avm_address        (cnn_top_0_load_read_avalon_address),                  //   load_read_avalon.address
		.load_avm_burstcount     (cnn_top_0_load_read_avalon_burstcount),               //                   .burstcount
		.load_avm_byteenable     (cnn_top_0_load_read_avalon_byteenable),               //                   .byteenable
		.load_avm_read           (cnn_top_0_load_read_avalon_read),                     //                   .read
		.load_avm_readdata       (cnn_top_0_load_read_avalon_readdata),                 //                   .readdata
		.load_avm_readdatavalid  (cnn_top_0_load_read_avalon_readdatavalid),            //                   .readdatavalid
		.load_avm_waitrequest    (cnn_top_0_load_read_avalon_waitrequest),              //                   .waitrequest
		.output_avm_address      (cnn_top_0_output_read_avalon_address),                // output_read_avalon.address
		.output_avm_burstcount   (cnn_top_0_output_read_avalon_burstcount),             //                   .burstcount
		.output_avm_byteenable   (cnn_top_0_output_read_avalon_byteenable),             //                   .byteenable
		.output_avm_waitrequest  (cnn_top_0_output_read_avalon_waitrequest),            //                   .waitrequest
		.output_avm_write        (cnn_top_0_output_read_avalon_write),                  //                   .write
		.output_avm_writedata    (cnn_top_0_output_read_avalon_writedata),              //                   .writedata
		.scale_avm_waitrequest   (cnn_top_0_scale_avm_avalon_waitrequest),              //   scale_avm_avalon.waitrequest
		.scale_avm_readdatavalid (cnn_top_0_scale_avm_avalon_readdatavalid),            //                   .readdatavalid
		.scale_avm_readdata      (cnn_top_0_scale_avm_avalon_readdata),                 //                   .readdata
		.scale_avm_address       (cnn_top_0_scale_avm_avalon_address),                  //                   .address
		.scale_avm_read          (cnn_top_0_scale_avm_avalon_read),                     //                   .read
		.scale_avm_byteenable    (cnn_top_0_scale_avm_avalon_byteenable),               //                   .byteenable
		.scale_avm_burstcount    (cnn_top_0_scale_avm_avalon_burstcount)                //                   .burstcount
	);

	ddr3_vga_top #(
		.BURST_LEN (16)
	) ddr3_vga_0 (
		.clk               (clk_50_clk),                                     //    clock.clk
		.avalon_write      (mm_interconnect_3_ddr3_vga_0_cfg_bus_write),     //  cfg_bus.write
		.avalon_read       (mm_interconnect_3_ddr3_vga_0_cfg_bus_read),      //         .read
		.avalon_addr       (mm_interconnect_3_ddr3_vga_0_cfg_bus_address),   //         .address
		.avalon_read_data  (mm_interconnect_3_ddr3_vga_0_cfg_bus_readdata),  //         .readdata
		.avalon_write_data (mm_interconnect_3_ddr3_vga_0_cfg_bus_writedata), //         .writedata
		.avl_waitrequest   (ddr3_vga_0_data_bus_waitrequest),                // data_bus.waitrequest
		.avl_addr          (ddr3_vga_0_data_bus_address),                    //         .address
		.avl_rdata_valid   (ddr3_vga_0_data_bus_readdatavalid),              //         .readdatavalid
		.avl_rdata         (ddr3_vga_0_data_bus_readdata),                   //         .readdata
		.avl_wdata         (ddr3_vga_0_data_bus_writedata),                  //         .writedata
		.avl_be            (ddr3_vga_0_data_bus_byteenable),                 //         .byteenable
		.avl_read_req      (ddr3_vga_0_data_bus_read),                       //         .read
		.avl_write_req     (ddr3_vga_0_data_bus_write),                      //         .write
		.avl_size          (ddr3_vga_0_data_bus_burstcount),                 //         .burstcount
		.vga_clk           (ddr3_vga_0_vga_bus_vga_clk),                     //  vga_bus.vga_clk
		.vga_de            (ddr3_vga_0_vga_bus_vga_de),                      //         .vga_de
		.vga_hsync         (ddr3_vga_0_vga_bus_vga_hsync),                   //         .vga_hsync
		.vga_rgb           (ddr3_vga_0_vga_bus_vga_rgb),                     //         .vga_rgb
		.vga_vsync         (ddr3_vga_0_vga_bus_vga_vsync),                   //         .vga_vsync
		.rst_n             (~rst_controller_reset_out_reset)                 //    reset.reset_n
	);

	soc_system_dipsw_pio dipsw_pio (
		.clk        (clk_50_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_3_dipsw_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_3_dipsw_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_3_dipsw_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_3_dipsw_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_3_dipsw_pio_s1_readdata),   //                    .readdata
		.out_port   (dipsw_pio_external_connection_export)       // external_connection.export
	);

	dvp_ddr3_top #(
		.BURST_LEN (16)
	) dvp_ddr3_0 (
		.clk               (clk_50_clk),                                     //    clock.clk
		.avalon_write      (mm_interconnect_3_dvp_ddr3_0_cfg_bus_write),     //  cfg_bus.write
		.avalon_read       (mm_interconnect_3_dvp_ddr3_0_cfg_bus_read),      //         .read
		.avalon_addr       (mm_interconnect_3_dvp_ddr3_0_cfg_bus_address),   //         .address
		.avalon_read_data  (mm_interconnect_3_dvp_ddr3_0_cfg_bus_readdata),  //         .readdata
		.avalon_write_data (mm_interconnect_3_dvp_ddr3_0_cfg_bus_writedata), //         .writedata
		.avl_waitrequest   (dvp_ddr3_0_data_bus_waitrequest),                // data_bus.waitrequest
		.avl_addr          (dvp_ddr3_0_data_bus_address),                    //         .address
		.avl_rdata_valid   (dvp_ddr3_0_data_bus_readdatavalid),              //         .readdatavalid
		.avl_rdata         (dvp_ddr3_0_data_bus_readdata),                   //         .readdata
		.avl_wdata         (dvp_ddr3_0_data_bus_writedata),                  //         .writedata
		.avl_be            (dvp_ddr3_0_data_bus_byteenable),                 //         .byteenable
		.avl_read_req      (dvp_ddr3_0_data_bus_read),                       //         .read
		.avl_write_req     (dvp_ddr3_0_data_bus_write),                      //         .write
		.avl_size          (dvp_ddr3_0_data_bus_burstcount),                 //         .burstcount
		.dvp_data          (vcam_0_dvp_bus_dvp_data),                        //  dvp_bus.dvp_data
		.dvp_href          (vcam_0_dvp_bus_dvp_href),                        //         .dvp_href
		.dvp_pclk          (vcam_0_dvp_bus_dvp_pclk),                        //         .dvp_pclk
		.dvp_vsync         (vcam_0_dvp_bus_dvp_vsync),                       //         .dvp_vsync
		.rst_n             (~rst_controller_reset_out_reset)                 //    reset.reset_n
	);

	soc_system_f2sdram_only_master #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) f2sdram_only_master (
		.clk_clk              (clk_50_clk),                               //          clk.clk
		.clk_reset_reset      (~reset_50_reset_n),                        //    clk_reset.reset
		.master_address       (f2sdram_only_master_master_address),       //       master.address
		.master_readdata      (f2sdram_only_master_master_readdata),      //             .readdata
		.master_read          (f2sdram_only_master_master_read),          //             .read
		.master_write         (f2sdram_only_master_master_write),         //             .write
		.master_writedata     (f2sdram_only_master_master_writedata),     //             .writedata
		.master_waitrequest   (f2sdram_only_master_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (f2sdram_only_master_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (f2sdram_only_master_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                          // master_reset.reset
	);

	soc_system_f2sdram_only_master #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) fpga_only_master (
		.clk_clk              (clk_50_clk),                            //          clk.clk
		.clk_reset_reset      (~reset_50_reset_n),                     //    clk_reset.reset
		.master_address       (fpga_only_master_master_address),       //       master.address
		.master_readdata      (fpga_only_master_master_readdata),      //             .readdata
		.master_read          (fpga_only_master_master_read),          //             .read
		.master_write         (fpga_only_master_master_write),         //             .write
		.master_writedata     (fpga_only_master_master_writedata),     //             .writedata
		.master_waitrequest   (fpga_only_master_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (fpga_only_master_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (fpga_only_master_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                       // master_reset.reset
	);

	soc_system_hps_0 #(
		.F2S_Width (3),
		.S2F_Width (3)
	) hps_0 (
		.h2f_loan_in               (hps_0_h2f_loan_io_in),                                  //         h2f_loan_io.in
		.h2f_loan_out              (hps_0_h2f_loan_io_out),                                 //                    .out
		.h2f_loan_oe               (hps_0_h2f_loan_io_oe),                                  //                    .oe
		.f2h_cold_rst_req_n        (hps_0_f2h_cold_reset_req_reset_n),                      //  f2h_cold_reset_req.reset_n
		.f2h_dbg_rst_req_n         (hps_0_f2h_debug_reset_req_reset_n),                     // f2h_debug_reset_req.reset_n
		.f2h_warm_rst_req_n        (hps_0_f2h_warm_reset_req_reset_n),                      //  f2h_warm_reset_req.reset_n
		.f2h_stm_hwevents          (hps_0_f2h_stm_hw_events_stm_hwevents),                  //   f2h_stm_hw_events.stm_hwevents
		.mem_a                     (memory_mem_a),                                          //              memory.mem_a
		.mem_ba                    (memory_mem_ba),                                         //                    .mem_ba
		.mem_ck                    (memory_mem_ck),                                         //                    .mem_ck
		.mem_ck_n                  (memory_mem_ck_n),                                       //                    .mem_ck_n
		.mem_cke                   (memory_mem_cke),                                        //                    .mem_cke
		.mem_cs_n                  (memory_mem_cs_n),                                       //                    .mem_cs_n
		.mem_ras_n                 (memory_mem_ras_n),                                      //                    .mem_ras_n
		.mem_cas_n                 (memory_mem_cas_n),                                      //                    .mem_cas_n
		.mem_we_n                  (memory_mem_we_n),                                       //                    .mem_we_n
		.mem_reset_n               (memory_mem_reset_n),                                    //                    .mem_reset_n
		.mem_dq                    (memory_mem_dq),                                         //                    .mem_dq
		.mem_dqs                   (memory_mem_dqs),                                        //                    .mem_dqs
		.mem_dqs_n                 (memory_mem_dqs_n),                                      //                    .mem_dqs_n
		.mem_odt                   (memory_mem_odt),                                        //                    .mem_odt
		.mem_dm                    (memory_mem_dm),                                         //                    .mem_dm
		.oct_rzqin                 (memory_oct_rzqin),                                      //                    .oct_rzqin
		.hps_io_emac1_inst_TX_CLK  (hps_0_hps_io_hps_io_emac1_inst_TX_CLK),                 //              hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0    (hps_0_hps_io_hps_io_emac1_inst_TXD0),                   //                    .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1    (hps_0_hps_io_hps_io_emac1_inst_TXD1),                   //                    .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2    (hps_0_hps_io_hps_io_emac1_inst_TXD2),                   //                    .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3    (hps_0_hps_io_hps_io_emac1_inst_TXD3),                   //                    .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0    (hps_0_hps_io_hps_io_emac1_inst_RXD0),                   //                    .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO    (hps_0_hps_io_hps_io_emac1_inst_MDIO),                   //                    .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC     (hps_0_hps_io_hps_io_emac1_inst_MDC),                    //                    .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL  (hps_0_hps_io_hps_io_emac1_inst_RX_CTL),                 //                    .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL  (hps_0_hps_io_hps_io_emac1_inst_TX_CTL),                 //                    .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK  (hps_0_hps_io_hps_io_emac1_inst_RX_CLK),                 //                    .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1    (hps_0_hps_io_hps_io_emac1_inst_RXD1),                   //                    .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2    (hps_0_hps_io_hps_io_emac1_inst_RXD2),                   //                    .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3    (hps_0_hps_io_hps_io_emac1_inst_RXD3),                   //                    .hps_io_emac1_inst_RXD3
		.hps_io_sdio_inst_CMD      (hps_0_hps_io_hps_io_sdio_inst_CMD),                     //                    .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0       (hps_0_hps_io_hps_io_sdio_inst_D0),                      //                    .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1       (hps_0_hps_io_hps_io_sdio_inst_D1),                      //                    .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK      (hps_0_hps_io_hps_io_sdio_inst_CLK),                     //                    .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2       (hps_0_hps_io_hps_io_sdio_inst_D2),                      //                    .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3       (hps_0_hps_io_hps_io_sdio_inst_D3),                      //                    .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0       (hps_0_hps_io_hps_io_usb1_inst_D0),                      //                    .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1       (hps_0_hps_io_hps_io_usb1_inst_D1),                      //                    .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2       (hps_0_hps_io_hps_io_usb1_inst_D2),                      //                    .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3       (hps_0_hps_io_hps_io_usb1_inst_D3),                      //                    .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4       (hps_0_hps_io_hps_io_usb1_inst_D4),                      //                    .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5       (hps_0_hps_io_hps_io_usb1_inst_D5),                      //                    .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6       (hps_0_hps_io_hps_io_usb1_inst_D6),                      //                    .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7       (hps_0_hps_io_hps_io_usb1_inst_D7),                      //                    .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK      (hps_0_hps_io_hps_io_usb1_inst_CLK),                     //                    .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP      (hps_0_hps_io_hps_io_usb1_inst_STP),                     //                    .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR      (hps_0_hps_io_hps_io_usb1_inst_DIR),                     //                    .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT      (hps_0_hps_io_hps_io_usb1_inst_NXT),                     //                    .hps_io_usb1_inst_NXT
		.hps_io_uart0_inst_RX      (hps_0_hps_io_hps_io_uart0_inst_RX),                     //                    .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX      (hps_0_hps_io_hps_io_uart0_inst_TX),                     //                    .hps_io_uart0_inst_TX
		.hps_io_gpio_inst_GPIO34   (hps_0_hps_io_hps_io_gpio_inst_GPIO34),                  //                    .hps_io_gpio_inst_GPIO34
		.hps_io_gpio_inst_GPIO35   (hps_0_hps_io_hps_io_gpio_inst_GPIO35),                  //                    .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO48   (hps_0_hps_io_hps_io_gpio_inst_GPIO48),                  //                    .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO51   (hps_0_hps_io_hps_io_gpio_inst_GPIO51),                  //                    .hps_io_gpio_inst_GPIO51
		.hps_io_gpio_inst_GPIO52   (hps_0_hps_io_hps_io_gpio_inst_GPIO52),                  //                    .hps_io_gpio_inst_GPIO52
		.hps_io_gpio_inst_GPIO53   (hps_0_hps_io_hps_io_gpio_inst_GPIO53),                  //                    .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54   (hps_0_hps_io_hps_io_gpio_inst_GPIO54),                  //                    .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_LOANIO00 (hps_0_hps_io_hps_io_gpio_inst_LOANIO00),                //                    .hps_io_gpio_inst_LOANIO00
		.hps_io_gpio_inst_LOANIO09 (hps_0_hps_io_hps_io_gpio_inst_LOANIO09),                //                    .hps_io_gpio_inst_LOANIO09
		.h2f_rst_n                 (hps_0_h2f_reset_reset_n),                               //           h2f_reset.reset_n
		.f2h_sdram0_clk            (clk_cnn_clk),                                           //    f2h_sdram0_clock.clk
		.f2h_sdram0_ADDRESS        (mm_interconnect_5_hps_0_f2h_sdram0_data_address),       //     f2h_sdram0_data.address
		.f2h_sdram0_BURSTCOUNT     (mm_interconnect_5_hps_0_f2h_sdram0_data_burstcount),    //                    .burstcount
		.f2h_sdram0_WAITREQUEST    (mm_interconnect_5_hps_0_f2h_sdram0_data_waitrequest),   //                    .waitrequest
		.f2h_sdram0_READDATA       (mm_interconnect_5_hps_0_f2h_sdram0_data_readdata),      //                    .readdata
		.f2h_sdram0_READDATAVALID  (mm_interconnect_5_hps_0_f2h_sdram0_data_readdatavalid), //                    .readdatavalid
		.f2h_sdram0_READ           (mm_interconnect_5_hps_0_f2h_sdram0_data_read),          //                    .read
		.f2h_sdram0_WRITEDATA      (mm_interconnect_5_hps_0_f2h_sdram0_data_writedata),     //                    .writedata
		.f2h_sdram0_BYTEENABLE     (mm_interconnect_5_hps_0_f2h_sdram0_data_byteenable),    //                    .byteenable
		.f2h_sdram0_WRITE          (mm_interconnect_5_hps_0_f2h_sdram0_data_write),         //                    .write
		.h2f_axi_clk               (clk_50_clk),                                            //       h2f_axi_clock.clk
		.h2f_AWID                  (),                                                      //      h2f_axi_master.awid
		.h2f_AWADDR                (),                                                      //                    .awaddr
		.h2f_AWLEN                 (),                                                      //                    .awlen
		.h2f_AWSIZE                (),                                                      //                    .awsize
		.h2f_AWBURST               (),                                                      //                    .awburst
		.h2f_AWLOCK                (),                                                      //                    .awlock
		.h2f_AWCACHE               (),                                                      //                    .awcache
		.h2f_AWPROT                (),                                                      //                    .awprot
		.h2f_AWVALID               (),                                                      //                    .awvalid
		.h2f_AWREADY               (),                                                      //                    .awready
		.h2f_WID                   (),                                                      //                    .wid
		.h2f_WDATA                 (),                                                      //                    .wdata
		.h2f_WSTRB                 (),                                                      //                    .wstrb
		.h2f_WLAST                 (),                                                      //                    .wlast
		.h2f_WVALID                (),                                                      //                    .wvalid
		.h2f_WREADY                (),                                                      //                    .wready
		.h2f_BID                   (),                                                      //                    .bid
		.h2f_BRESP                 (),                                                      //                    .bresp
		.h2f_BVALID                (),                                                      //                    .bvalid
		.h2f_BREADY                (),                                                      //                    .bready
		.h2f_ARID                  (),                                                      //                    .arid
		.h2f_ARADDR                (),                                                      //                    .araddr
		.h2f_ARLEN                 (),                                                      //                    .arlen
		.h2f_ARSIZE                (),                                                      //                    .arsize
		.h2f_ARBURST               (),                                                      //                    .arburst
		.h2f_ARLOCK                (),                                                      //                    .arlock
		.h2f_ARCACHE               (),                                                      //                    .arcache
		.h2f_ARPROT                (),                                                      //                    .arprot
		.h2f_ARVALID               (),                                                      //                    .arvalid
		.h2f_ARREADY               (),                                                      //                    .arready
		.h2f_RID                   (),                                                      //                    .rid
		.h2f_RDATA                 (),                                                      //                    .rdata
		.h2f_RRESP                 (),                                                      //                    .rresp
		.h2f_RLAST                 (),                                                      //                    .rlast
		.h2f_RVALID                (),                                                      //                    .rvalid
		.h2f_RREADY                (),                                                      //                    .rready
		.f2h_axi_clk               (clk_50_clk),                                            //       f2h_axi_clock.clk
		.f2h_AWID                  (mm_interconnect_4_hps_0_f2h_axi_slave_awid),            //       f2h_axi_slave.awid
		.f2h_AWADDR                (mm_interconnect_4_hps_0_f2h_axi_slave_awaddr),          //                    .awaddr
		.f2h_AWLEN                 (mm_interconnect_4_hps_0_f2h_axi_slave_awlen),           //                    .awlen
		.f2h_AWSIZE                (mm_interconnect_4_hps_0_f2h_axi_slave_awsize),          //                    .awsize
		.f2h_AWBURST               (mm_interconnect_4_hps_0_f2h_axi_slave_awburst),         //                    .awburst
		.f2h_AWLOCK                (mm_interconnect_4_hps_0_f2h_axi_slave_awlock),          //                    .awlock
		.f2h_AWCACHE               (mm_interconnect_4_hps_0_f2h_axi_slave_awcache),         //                    .awcache
		.f2h_AWPROT                (mm_interconnect_4_hps_0_f2h_axi_slave_awprot),          //                    .awprot
		.f2h_AWVALID               (mm_interconnect_4_hps_0_f2h_axi_slave_awvalid),         //                    .awvalid
		.f2h_AWREADY               (mm_interconnect_4_hps_0_f2h_axi_slave_awready),         //                    .awready
		.f2h_AWUSER                (mm_interconnect_4_hps_0_f2h_axi_slave_awuser),          //                    .awuser
		.f2h_WID                   (mm_interconnect_4_hps_0_f2h_axi_slave_wid),             //                    .wid
		.f2h_WDATA                 (mm_interconnect_4_hps_0_f2h_axi_slave_wdata),           //                    .wdata
		.f2h_WSTRB                 (mm_interconnect_4_hps_0_f2h_axi_slave_wstrb),           //                    .wstrb
		.f2h_WLAST                 (mm_interconnect_4_hps_0_f2h_axi_slave_wlast),           //                    .wlast
		.f2h_WVALID                (mm_interconnect_4_hps_0_f2h_axi_slave_wvalid),          //                    .wvalid
		.f2h_WREADY                (mm_interconnect_4_hps_0_f2h_axi_slave_wready),          //                    .wready
		.f2h_BID                   (mm_interconnect_4_hps_0_f2h_axi_slave_bid),             //                    .bid
		.f2h_BRESP                 (mm_interconnect_4_hps_0_f2h_axi_slave_bresp),           //                    .bresp
		.f2h_BVALID                (mm_interconnect_4_hps_0_f2h_axi_slave_bvalid),          //                    .bvalid
		.f2h_BREADY                (mm_interconnect_4_hps_0_f2h_axi_slave_bready),          //                    .bready
		.f2h_ARID                  (mm_interconnect_4_hps_0_f2h_axi_slave_arid),            //                    .arid
		.f2h_ARADDR                (mm_interconnect_4_hps_0_f2h_axi_slave_araddr),          //                    .araddr
		.f2h_ARLEN                 (mm_interconnect_4_hps_0_f2h_axi_slave_arlen),           //                    .arlen
		.f2h_ARSIZE                (mm_interconnect_4_hps_0_f2h_axi_slave_arsize),          //                    .arsize
		.f2h_ARBURST               (mm_interconnect_4_hps_0_f2h_axi_slave_arburst),         //                    .arburst
		.f2h_ARLOCK                (mm_interconnect_4_hps_0_f2h_axi_slave_arlock),          //                    .arlock
		.f2h_ARCACHE               (mm_interconnect_4_hps_0_f2h_axi_slave_arcache),         //                    .arcache
		.f2h_ARPROT                (mm_interconnect_4_hps_0_f2h_axi_slave_arprot),          //                    .arprot
		.f2h_ARVALID               (mm_interconnect_4_hps_0_f2h_axi_slave_arvalid),         //                    .arvalid
		.f2h_ARREADY               (mm_interconnect_4_hps_0_f2h_axi_slave_arready),         //                    .arready
		.f2h_ARUSER                (mm_interconnect_4_hps_0_f2h_axi_slave_aruser),          //                    .aruser
		.f2h_RID                   (mm_interconnect_4_hps_0_f2h_axi_slave_rid),             //                    .rid
		.f2h_RDATA                 (mm_interconnect_4_hps_0_f2h_axi_slave_rdata),           //                    .rdata
		.f2h_RRESP                 (mm_interconnect_4_hps_0_f2h_axi_slave_rresp),           //                    .rresp
		.f2h_RLAST                 (mm_interconnect_4_hps_0_f2h_axi_slave_rlast),           //                    .rlast
		.f2h_RVALID                (mm_interconnect_4_hps_0_f2h_axi_slave_rvalid),          //                    .rvalid
		.f2h_RREADY                (mm_interconnect_4_hps_0_f2h_axi_slave_rready),          //                    .rready
		.h2f_lw_axi_clk            (clk_50_clk),                                            //    h2f_lw_axi_clock.clk
		.h2f_lw_AWID               (hps_0_h2f_lw_axi_master_awid),                          //   h2f_lw_axi_master.awid
		.h2f_lw_AWADDR             (hps_0_h2f_lw_axi_master_awaddr),                        //                    .awaddr
		.h2f_lw_AWLEN              (hps_0_h2f_lw_axi_master_awlen),                         //                    .awlen
		.h2f_lw_AWSIZE             (hps_0_h2f_lw_axi_master_awsize),                        //                    .awsize
		.h2f_lw_AWBURST            (hps_0_h2f_lw_axi_master_awburst),                       //                    .awburst
		.h2f_lw_AWLOCK             (hps_0_h2f_lw_axi_master_awlock),                        //                    .awlock
		.h2f_lw_AWCACHE            (hps_0_h2f_lw_axi_master_awcache),                       //                    .awcache
		.h2f_lw_AWPROT             (hps_0_h2f_lw_axi_master_awprot),                        //                    .awprot
		.h2f_lw_AWVALID            (hps_0_h2f_lw_axi_master_awvalid),                       //                    .awvalid
		.h2f_lw_AWREADY            (hps_0_h2f_lw_axi_master_awready),                       //                    .awready
		.h2f_lw_WID                (hps_0_h2f_lw_axi_master_wid),                           //                    .wid
		.h2f_lw_WDATA              (hps_0_h2f_lw_axi_master_wdata),                         //                    .wdata
		.h2f_lw_WSTRB              (hps_0_h2f_lw_axi_master_wstrb),                         //                    .wstrb
		.h2f_lw_WLAST              (hps_0_h2f_lw_axi_master_wlast),                         //                    .wlast
		.h2f_lw_WVALID             (hps_0_h2f_lw_axi_master_wvalid),                        //                    .wvalid
		.h2f_lw_WREADY             (hps_0_h2f_lw_axi_master_wready),                        //                    .wready
		.h2f_lw_BID                (hps_0_h2f_lw_axi_master_bid),                           //                    .bid
		.h2f_lw_BRESP              (hps_0_h2f_lw_axi_master_bresp),                         //                    .bresp
		.h2f_lw_BVALID             (hps_0_h2f_lw_axi_master_bvalid),                        //                    .bvalid
		.h2f_lw_BREADY             (hps_0_h2f_lw_axi_master_bready),                        //                    .bready
		.h2f_lw_ARID               (hps_0_h2f_lw_axi_master_arid),                          //                    .arid
		.h2f_lw_ARADDR             (hps_0_h2f_lw_axi_master_araddr),                        //                    .araddr
		.h2f_lw_ARLEN              (hps_0_h2f_lw_axi_master_arlen),                         //                    .arlen
		.h2f_lw_ARSIZE             (hps_0_h2f_lw_axi_master_arsize),                        //                    .arsize
		.h2f_lw_ARBURST            (hps_0_h2f_lw_axi_master_arburst),                       //                    .arburst
		.h2f_lw_ARLOCK             (hps_0_h2f_lw_axi_master_arlock),                        //                    .arlock
		.h2f_lw_ARCACHE            (hps_0_h2f_lw_axi_master_arcache),                       //                    .arcache
		.h2f_lw_ARPROT             (hps_0_h2f_lw_axi_master_arprot),                        //                    .arprot
		.h2f_lw_ARVALID            (hps_0_h2f_lw_axi_master_arvalid),                       //                    .arvalid
		.h2f_lw_ARREADY            (hps_0_h2f_lw_axi_master_arready),                       //                    .arready
		.h2f_lw_RID                (hps_0_h2f_lw_axi_master_rid),                           //                    .rid
		.h2f_lw_RDATA              (hps_0_h2f_lw_axi_master_rdata),                         //                    .rdata
		.h2f_lw_RRESP              (hps_0_h2f_lw_axi_master_rresp),                         //                    .rresp
		.h2f_lw_RLAST              (hps_0_h2f_lw_axi_master_rlast),                         //                    .rlast
		.h2f_lw_RVALID             (hps_0_h2f_lw_axi_master_rvalid),                        //                    .rvalid
		.h2f_lw_RREADY             (hps_0_h2f_lw_axi_master_rready),                        //                    .rready
		.f2h_irq_p0                (hps_0_f2h_irq0_irq),                                    //            f2h_irq0.irq
		.f2h_irq_p1                (hps_0_f2h_irq1_irq)                                     //            f2h_irq1.irq
	);

	soc_system_f2sdram_only_master #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) hps_only_master (
		.clk_clk              (clk_50_clk),                           //          clk.clk
		.clk_reset_reset      (~reset_50_reset_n),                    //    clk_reset.reset
		.master_address       (hps_only_master_master_address),       //       master.address
		.master_readdata      (hps_only_master_master_readdata),      //             .readdata
		.master_read          (hps_only_master_master_read),          //             .read
		.master_write         (hps_only_master_master_write),         //             .write
		.master_writedata     (hps_only_master_master_writedata),     //             .writedata
		.master_waitrequest   (hps_only_master_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (hps_only_master_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (hps_only_master_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                      // master_reset.reset
	);

	soc_system_led_pio led_pio (
		.clk        (clk_50_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_3_led_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_3_led_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_3_led_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_3_led_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_3_led_pio_s1_readdata),   //                    .readdata
		.in_port    (led_pio_external_connection_export)       // external_connection.export
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (128),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (32),
		.BURSTCOUNT_WIDTH  (5),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_axi (
		.clk              (clk_50_clk),                                       //   clk.clk
		.reset            (rst_controller_reset_out_reset),                   // reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_bridge_axi_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_bridge_axi_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_bridge_axi_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_bridge_axi_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_mm_bridge_axi_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_mm_bridge_axi_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_mm_bridge_axi_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_mm_bridge_axi_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_mm_bridge_axi_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_bridge_axi_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mm_bridge_axi_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (mm_bridge_axi_m0_readdata),                        //      .readdata
		.m0_readdatavalid (mm_bridge_axi_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (mm_bridge_axi_m0_burstcount),                      //      .burstcount
		.m0_writedata     (mm_bridge_axi_m0_writedata),                       //      .writedata
		.m0_address       (mm_bridge_axi_m0_address),                         //      .address
		.m0_write         (mm_bridge_axi_m0_write),                           //      .write
		.m0_read          (mm_bridge_axi_m0_read),                            //      .read
		.m0_byteenable    (mm_bridge_axi_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (mm_bridge_axi_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                                 // (terminated)
		.m0_response      (2'b00)                                             // (terminated)
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (15),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_lw_axi (
		.clk              (clk_50_clk),                                          //   clk.clk
		.reset            (rst_controller_reset_out_reset),                      // reset.reset
		.s0_waitrequest   (mm_interconnect_1_mm_bridge_lw_axi_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_1_mm_bridge_lw_axi_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_1_mm_bridge_lw_axi_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_1_mm_bridge_lw_axi_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_1_mm_bridge_lw_axi_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_1_mm_bridge_lw_axi_s0_address),       //      .address
		.s0_write         (mm_interconnect_1_mm_bridge_lw_axi_s0_write),         //      .write
		.s0_read          (mm_interconnect_1_mm_bridge_lw_axi_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_1_mm_bridge_lw_axi_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_1_mm_bridge_lw_axi_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mm_bridge_lw_axi_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (mm_bridge_lw_axi_m0_readdata),                        //      .readdata
		.m0_readdatavalid (mm_bridge_lw_axi_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (mm_bridge_lw_axi_m0_burstcount),                      //      .burstcount
		.m0_writedata     (mm_bridge_lw_axi_m0_writedata),                       //      .writedata
		.m0_address       (mm_bridge_lw_axi_m0_address),                         //      .address
		.m0_write         (mm_bridge_lw_axi_m0_write),                           //      .write
		.m0_read          (mm_bridge_lw_axi_m0_read),                            //      .read
		.m0_byteenable    (mm_bridge_lw_axi_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (mm_bridge_lw_axi_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                                    // (terminated)
		.m0_response      (2'b00)                                                // (terminated)
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (128),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (32),
		.BURSTCOUNT_WIDTH  (5),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_sdram0 (
		.clk              (clk_cnn_clk),                                         //   clk.clk
		.reset            (rst_controller_001_reset_out_reset),                  // reset.reset
		.s0_waitrequest   (mm_interconnect_2_mm_bridge_sdram0_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_2_mm_bridge_sdram0_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_2_mm_bridge_sdram0_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_2_mm_bridge_sdram0_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_2_mm_bridge_sdram0_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_2_mm_bridge_sdram0_s0_address),       //      .address
		.s0_write         (mm_interconnect_2_mm_bridge_sdram0_s0_write),         //      .write
		.s0_read          (mm_interconnect_2_mm_bridge_sdram0_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_2_mm_bridge_sdram0_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_2_mm_bridge_sdram0_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mm_bridge_sdram0_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (mm_bridge_sdram0_m0_readdata),                        //      .readdata
		.m0_readdatavalid (mm_bridge_sdram0_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (mm_bridge_sdram0_m0_burstcount),                      //      .burstcount
		.m0_writedata     (mm_bridge_sdram0_m0_writedata),                       //      .writedata
		.m0_address       (mm_bridge_sdram0_m0_address),                         //      .address
		.m0_write         (mm_bridge_sdram0_m0_write),                           //      .write
		.m0_read          (mm_bridge_sdram0_m0_read),                            //      .read
		.m0_byteenable    (mm_bridge_sdram0_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (mm_bridge_sdram0_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                                    // (terminated)
		.m0_response      (2'b00)                                                // (terminated)
	);

	soc_system_sld_hub_controller_system_0 #(
		.ENABLE_JTAG_IO_SELECTION (0)
	) sld_hub_controller_system_0 (
		.clk_clk          (clk_50_clk),                                                     //   clk.clk
		.reset_reset      (rst_controller_reset_out_reset),                                 // reset.reset
		.s0_waitrequest   (mm_interconnect_3_sld_hub_controller_system_0_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_3_sld_hub_controller_system_0_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_3_sld_hub_controller_system_0_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_3_sld_hub_controller_system_0_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_3_sld_hub_controller_system_0_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_3_sld_hub_controller_system_0_s0_address),       //      .address
		.s0_write         (mm_interconnect_3_sld_hub_controller_system_0_s0_write),         //      .write
		.s0_read          (mm_interconnect_3_sld_hub_controller_system_0_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_3_sld_hub_controller_system_0_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_3_sld_hub_controller_system_0_s0_debugaccess)    //      .debugaccess
	);

	soc_system_sysid_qsys sysid_qsys (
		.clock    (clk_50_clk),                                          //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.readdata (mm_interconnect_3_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_3_sysid_qsys_control_slave_address)   //              .address
	);

	vcam_top #(
		.BURST_LEN (16)
	) vcam_0 (
		.clk             (clk_50_clk),                                 //    clock.clk
		.avm_write       (vcam_0_data_bus_write),                      // data_bus.write
		.avm_read        (vcam_0_data_bus_read),                       //         .read
		.avm_addr        (vcam_0_data_bus_address),                    //         .address
		.avm_waitrequest (vcam_0_data_bus_waitrequest),                //         .waitrequest
		.avm_rdata_valid (vcam_0_data_bus_readdatavalid),              //         .readdatavalid
		.avm_rdata       (vcam_0_data_bus_readdata),                   //         .readdata
		.avm_wdata       (vcam_0_data_bus_writedata),                  //         .writedata
		.avm_byteenable  (vcam_0_data_bus_byteenable),                 //         .byteenable
		.avm_size        (vcam_0_data_bus_burstcount),                 //         .burstcount
		.cfg_addr        (mm_interconnect_3_vcam_0_cfg_bus_address),   //  cfg_bus.address
		.cfg_write_data  (mm_interconnect_3_vcam_0_cfg_bus_writedata), //         .writedata
		.cfg_read_data   (mm_interconnect_3_vcam_0_cfg_bus_readdata),  //         .readdata
		.cfg_read        (mm_interconnect_3_vcam_0_cfg_bus_read),      //         .read
		.cfg_write       (mm_interconnect_3_vcam_0_cfg_bus_write),     //         .write
		.dvp_data        (vcam_0_dvp_bus_dvp_data),                    //  dvp_bus.dvp_data
		.dvp_href        (vcam_0_dvp_bus_dvp_href),                    //         .dvp_href
		.dvp_pclk        (vcam_0_dvp_bus_dvp_pclk),                    //         .dvp_pclk
		.dvp_vsync       (vcam_0_dvp_bus_dvp_vsync),                   //         .dvp_vsync
		.rst_n           (~rst_controller_reset_out_reset)             //    reset.reset_n
	);

	receive_top #(
		.BUF1_BASE_ADDR (0),
		.BUF2_BASE_ADDR (384000)
	) vhdmi_0 (
		.s_avl_wr_req      (mm_interconnect_3_vhdmi_0_s_avalon_mm_write),      // s_avalon_mm.write
		.s_avl_rd_req      (mm_interconnect_3_vhdmi_0_s_avalon_mm_read),       //            .read
		.s_avl_wr_data     (mm_interconnect_3_vhdmi_0_s_avalon_mm_writedata),  //            .writedata
		.s_avl_rd_data     (mm_interconnect_3_vhdmi_0_s_avalon_mm_readdata),   //            .readdata
		.s_avl_address     (mm_interconnect_3_vhdmi_0_s_avalon_mm_address),    //            .address
		.s_avl_chipselect  (mm_interconnect_3_vhdmi_0_s_avalon_mm_chipselect), //            .chipselect
		.m_avl_addr        (vhdmi_0_m_avalon_mm_address),                      // m_avalon_mm.address
		.m_avl_be          (vhdmi_0_m_avalon_mm_byteenable),                   //            .byteenable
		.m_avl_size        (vhdmi_0_m_avalon_mm_burstcount),                   //            .burstcount
		.m_avl_wdata       (vhdmi_0_m_avalon_mm_writedata),                    //            .writedata
		.m_avl_write_req   (vhdmi_0_m_avalon_mm_write),                        //            .write
		.m_avl_waitrequest (vhdmi_0_m_avalon_mm_waitrequest),                  //            .waitrequest
		.rst_n             (~rst_controller_reset_out_reset),                  //       rst_n.reset_n
		.vga_clk           (ddr3_vga_0_vga_bus_vga_clk),                       //      vga_in.vga_clk
		.vga_de            (ddr3_vga_0_vga_bus_vga_de),                        //            .vga_de
		.vga_hsync         (ddr3_vga_0_vga_bus_vga_hsync),                     //            .vga_hsync
		.vga_vsync         (ddr3_vga_0_vga_bus_vga_vsync),                     //            .vga_vsync
		.vga_rgb           (ddr3_vga_0_vga_bus_vga_rgb),                       //            .vga_rgb
		.clk_hps           (clk_50_clk)                                        //     clk_hps.clk
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_50_clk_clk                           (clk_50_clk),                                       //                         clk_50_clk.clk
		.vcam_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                   // vcam_0_reset_reset_bridge_in_reset.reset
		.ddr3_vga_0_data_bus_address              (ddr3_vga_0_data_bus_address),                      //                ddr3_vga_0_data_bus.address
		.ddr3_vga_0_data_bus_waitrequest          (ddr3_vga_0_data_bus_waitrequest),                  //                                   .waitrequest
		.ddr3_vga_0_data_bus_burstcount           (ddr3_vga_0_data_bus_burstcount),                   //                                   .burstcount
		.ddr3_vga_0_data_bus_byteenable           (ddr3_vga_0_data_bus_byteenable),                   //                                   .byteenable
		.ddr3_vga_0_data_bus_read                 (ddr3_vga_0_data_bus_read),                         //                                   .read
		.ddr3_vga_0_data_bus_readdata             (ddr3_vga_0_data_bus_readdata),                     //                                   .readdata
		.ddr3_vga_0_data_bus_readdatavalid        (ddr3_vga_0_data_bus_readdatavalid),                //                                   .readdatavalid
		.ddr3_vga_0_data_bus_write                (ddr3_vga_0_data_bus_write),                        //                                   .write
		.ddr3_vga_0_data_bus_writedata            (ddr3_vga_0_data_bus_writedata),                    //                                   .writedata
		.dvp_ddr3_0_data_bus_address              (dvp_ddr3_0_data_bus_address),                      //                dvp_ddr3_0_data_bus.address
		.dvp_ddr3_0_data_bus_waitrequest          (dvp_ddr3_0_data_bus_waitrequest),                  //                                   .waitrequest
		.dvp_ddr3_0_data_bus_burstcount           (dvp_ddr3_0_data_bus_burstcount),                   //                                   .burstcount
		.dvp_ddr3_0_data_bus_byteenable           (dvp_ddr3_0_data_bus_byteenable),                   //                                   .byteenable
		.dvp_ddr3_0_data_bus_read                 (dvp_ddr3_0_data_bus_read),                         //                                   .read
		.dvp_ddr3_0_data_bus_readdata             (dvp_ddr3_0_data_bus_readdata),                     //                                   .readdata
		.dvp_ddr3_0_data_bus_readdatavalid        (dvp_ddr3_0_data_bus_readdatavalid),                //                                   .readdatavalid
		.dvp_ddr3_0_data_bus_write                (dvp_ddr3_0_data_bus_write),                        //                                   .write
		.dvp_ddr3_0_data_bus_writedata            (dvp_ddr3_0_data_bus_writedata),                    //                                   .writedata
		.vcam_0_data_bus_address                  (vcam_0_data_bus_address),                          //                    vcam_0_data_bus.address
		.vcam_0_data_bus_waitrequest              (vcam_0_data_bus_waitrequest),                      //                                   .waitrequest
		.vcam_0_data_bus_burstcount               (vcam_0_data_bus_burstcount),                       //                                   .burstcount
		.vcam_0_data_bus_byteenable               (vcam_0_data_bus_byteenable),                       //                                   .byteenable
		.vcam_0_data_bus_read                     (vcam_0_data_bus_read),                             //                                   .read
		.vcam_0_data_bus_readdata                 (vcam_0_data_bus_readdata),                         //                                   .readdata
		.vcam_0_data_bus_readdatavalid            (vcam_0_data_bus_readdatavalid),                    //                                   .readdatavalid
		.vcam_0_data_bus_write                    (vcam_0_data_bus_write),                            //                                   .write
		.vcam_0_data_bus_writedata                (vcam_0_data_bus_writedata),                        //                                   .writedata
		.vhdmi_0_m_avalon_mm_address              (vhdmi_0_m_avalon_mm_address),                      //                vhdmi_0_m_avalon_mm.address
		.vhdmi_0_m_avalon_mm_waitrequest          (vhdmi_0_m_avalon_mm_waitrequest),                  //                                   .waitrequest
		.vhdmi_0_m_avalon_mm_burstcount           (vhdmi_0_m_avalon_mm_burstcount),                   //                                   .burstcount
		.vhdmi_0_m_avalon_mm_byteenable           (vhdmi_0_m_avalon_mm_byteenable),                   //                                   .byteenable
		.vhdmi_0_m_avalon_mm_write                (vhdmi_0_m_avalon_mm_write),                        //                                   .write
		.vhdmi_0_m_avalon_mm_writedata            (vhdmi_0_m_avalon_mm_writedata),                    //                                   .writedata
		.mm_bridge_axi_s0_address                 (mm_interconnect_0_mm_bridge_axi_s0_address),       //                   mm_bridge_axi_s0.address
		.mm_bridge_axi_s0_write                   (mm_interconnect_0_mm_bridge_axi_s0_write),         //                                   .write
		.mm_bridge_axi_s0_read                    (mm_interconnect_0_mm_bridge_axi_s0_read),          //                                   .read
		.mm_bridge_axi_s0_readdata                (mm_interconnect_0_mm_bridge_axi_s0_readdata),      //                                   .readdata
		.mm_bridge_axi_s0_writedata               (mm_interconnect_0_mm_bridge_axi_s0_writedata),     //                                   .writedata
		.mm_bridge_axi_s0_burstcount              (mm_interconnect_0_mm_bridge_axi_s0_burstcount),    //                                   .burstcount
		.mm_bridge_axi_s0_byteenable              (mm_interconnect_0_mm_bridge_axi_s0_byteenable),    //                                   .byteenable
		.mm_bridge_axi_s0_readdatavalid           (mm_interconnect_0_mm_bridge_axi_s0_readdatavalid), //                                   .readdatavalid
		.mm_bridge_axi_s0_waitrequest             (mm_interconnect_0_mm_bridge_axi_s0_waitrequest),   //                                   .waitrequest
		.mm_bridge_axi_s0_debugaccess             (mm_interconnect_0_mm_bridge_axi_s0_debugaccess)    //                                   .debugaccess
	);

	soc_system_mm_interconnect_1 mm_interconnect_1 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                        //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                      //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                       //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                      //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                     //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                      //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                     //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                      //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                     //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                     //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                         //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                       //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                       //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                       //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                      //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                      //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                         //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                       //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                      //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                      //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                        //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                      //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                       //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                      //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                     //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                      //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                     //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                      //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                     //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                     //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                         //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                       //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                       //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                       //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                      //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                      //                                                              .rready
		.clk_50_clk_clk                                                      (clk_50_clk),                                          //                                                    clk_50_clk.clk
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                  // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.mm_bridge_lw_axi_reset_reset_bridge_in_reset_reset                  (rst_controller_reset_out_reset),                      //                  mm_bridge_lw_axi_reset_reset_bridge_in_reset.reset
		.mm_bridge_lw_axi_s0_address                                         (mm_interconnect_1_mm_bridge_lw_axi_s0_address),       //                                           mm_bridge_lw_axi_s0.address
		.mm_bridge_lw_axi_s0_write                                           (mm_interconnect_1_mm_bridge_lw_axi_s0_write),         //                                                              .write
		.mm_bridge_lw_axi_s0_read                                            (mm_interconnect_1_mm_bridge_lw_axi_s0_read),          //                                                              .read
		.mm_bridge_lw_axi_s0_readdata                                        (mm_interconnect_1_mm_bridge_lw_axi_s0_readdata),      //                                                              .readdata
		.mm_bridge_lw_axi_s0_writedata                                       (mm_interconnect_1_mm_bridge_lw_axi_s0_writedata),     //                                                              .writedata
		.mm_bridge_lw_axi_s0_burstcount                                      (mm_interconnect_1_mm_bridge_lw_axi_s0_burstcount),    //                                                              .burstcount
		.mm_bridge_lw_axi_s0_byteenable                                      (mm_interconnect_1_mm_bridge_lw_axi_s0_byteenable),    //                                                              .byteenable
		.mm_bridge_lw_axi_s0_readdatavalid                                   (mm_interconnect_1_mm_bridge_lw_axi_s0_readdatavalid), //                                                              .readdatavalid
		.mm_bridge_lw_axi_s0_waitrequest                                     (mm_interconnect_1_mm_bridge_lw_axi_s0_waitrequest),   //                                                              .waitrequest
		.mm_bridge_lw_axi_s0_debugaccess                                     (mm_interconnect_1_mm_bridge_lw_axi_s0_debugaccess)    //                                                              .debugaccess
	);

	soc_system_mm_interconnect_2 mm_interconnect_2 (
		.clk_cnn_clk_clk                             (clk_cnn_clk),                                         //                           clk_cnn_clk.clk
		.cnn_top_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                  // cnn_top_0_reset_reset_bridge_in_reset.reset
		.cnn_top_0_load_read_avalon_address          (cnn_top_0_load_read_avalon_address),                  //            cnn_top_0_load_read_avalon.address
		.cnn_top_0_load_read_avalon_waitrequest      (cnn_top_0_load_read_avalon_waitrequest),              //                                      .waitrequest
		.cnn_top_0_load_read_avalon_burstcount       (cnn_top_0_load_read_avalon_burstcount),               //                                      .burstcount
		.cnn_top_0_load_read_avalon_byteenable       (cnn_top_0_load_read_avalon_byteenable),               //                                      .byteenable
		.cnn_top_0_load_read_avalon_read             (cnn_top_0_load_read_avalon_read),                     //                                      .read
		.cnn_top_0_load_read_avalon_readdata         (cnn_top_0_load_read_avalon_readdata),                 //                                      .readdata
		.cnn_top_0_load_read_avalon_readdatavalid    (cnn_top_0_load_read_avalon_readdatavalid),            //                                      .readdatavalid
		.cnn_top_0_output_read_avalon_address        (cnn_top_0_output_read_avalon_address),                //          cnn_top_0_output_read_avalon.address
		.cnn_top_0_output_read_avalon_waitrequest    (cnn_top_0_output_read_avalon_waitrequest),            //                                      .waitrequest
		.cnn_top_0_output_read_avalon_burstcount     (cnn_top_0_output_read_avalon_burstcount),             //                                      .burstcount
		.cnn_top_0_output_read_avalon_byteenable     (cnn_top_0_output_read_avalon_byteenable),             //                                      .byteenable
		.cnn_top_0_output_read_avalon_write          (cnn_top_0_output_read_avalon_write),                  //                                      .write
		.cnn_top_0_output_read_avalon_writedata      (cnn_top_0_output_read_avalon_writedata),              //                                      .writedata
		.cnn_top_0_param_read_avalon_address         (cnn_top_0_param_read_avalon_address),                 //           cnn_top_0_param_read_avalon.address
		.cnn_top_0_param_read_avalon_waitrequest     (cnn_top_0_param_read_avalon_waitrequest),             //                                      .waitrequest
		.cnn_top_0_param_read_avalon_burstcount      (cnn_top_0_param_read_avalon_burstcount),              //                                      .burstcount
		.cnn_top_0_param_read_avalon_byteenable      (cnn_top_0_param_read_avalon_byteenable),              //                                      .byteenable
		.cnn_top_0_param_read_avalon_read            (cnn_top_0_param_read_avalon_read),                    //                                      .read
		.cnn_top_0_param_read_avalon_readdata        (cnn_top_0_param_read_avalon_readdata),                //                                      .readdata
		.cnn_top_0_param_read_avalon_readdatavalid   (cnn_top_0_param_read_avalon_readdatavalid),           //                                      .readdatavalid
		.cnn_top_0_scale_avm_avalon_address          (cnn_top_0_scale_avm_avalon_address),                  //            cnn_top_0_scale_avm_avalon.address
		.cnn_top_0_scale_avm_avalon_waitrequest      (cnn_top_0_scale_avm_avalon_waitrequest),              //                                      .waitrequest
		.cnn_top_0_scale_avm_avalon_burstcount       (cnn_top_0_scale_avm_avalon_burstcount),               //                                      .burstcount
		.cnn_top_0_scale_avm_avalon_byteenable       (cnn_top_0_scale_avm_avalon_byteenable),               //                                      .byteenable
		.cnn_top_0_scale_avm_avalon_read             (cnn_top_0_scale_avm_avalon_read),                     //                                      .read
		.cnn_top_0_scale_avm_avalon_readdata         (cnn_top_0_scale_avm_avalon_readdata),                 //                                      .readdata
		.cnn_top_0_scale_avm_avalon_readdatavalid    (cnn_top_0_scale_avm_avalon_readdatavalid),            //                                      .readdatavalid
		.mm_bridge_sdram0_s0_address                 (mm_interconnect_2_mm_bridge_sdram0_s0_address),       //                   mm_bridge_sdram0_s0.address
		.mm_bridge_sdram0_s0_write                   (mm_interconnect_2_mm_bridge_sdram0_s0_write),         //                                      .write
		.mm_bridge_sdram0_s0_read                    (mm_interconnect_2_mm_bridge_sdram0_s0_read),          //                                      .read
		.mm_bridge_sdram0_s0_readdata                (mm_interconnect_2_mm_bridge_sdram0_s0_readdata),      //                                      .readdata
		.mm_bridge_sdram0_s0_writedata               (mm_interconnect_2_mm_bridge_sdram0_s0_writedata),     //                                      .writedata
		.mm_bridge_sdram0_s0_burstcount              (mm_interconnect_2_mm_bridge_sdram0_s0_burstcount),    //                                      .burstcount
		.mm_bridge_sdram0_s0_byteenable              (mm_interconnect_2_mm_bridge_sdram0_s0_byteenable),    //                                      .byteenable
		.mm_bridge_sdram0_s0_readdatavalid           (mm_interconnect_2_mm_bridge_sdram0_s0_readdatavalid), //                                      .readdatavalid
		.mm_bridge_sdram0_s0_waitrequest             (mm_interconnect_2_mm_bridge_sdram0_s0_waitrequest),   //                                      .waitrequest
		.mm_bridge_sdram0_s0_debugaccess             (mm_interconnect_2_mm_bridge_sdram0_s0_debugaccess)    //                                      .debugaccess
	);

	soc_system_mm_interconnect_3 mm_interconnect_3 (
		.clk_50_clk_clk                                         (clk_50_clk),                                                     //                                       clk_50_clk.clk
		.clk_cnn_clk_clk                                        (clk_cnn_clk),                                                    //                                      clk_cnn_clk.clk
		.cnn_top_0_reset_reset_bridge_in_reset_reset            (rst_controller_001_reset_out_reset),                             //            cnn_top_0_reset_reset_bridge_in_reset.reset
		.fpga_only_master_clk_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                 // fpga_only_master_clk_reset_reset_bridge_in_reset.reset
		.mm_bridge_lw_axi_reset_reset_bridge_in_reset_reset     (rst_controller_reset_out_reset),                                 //     mm_bridge_lw_axi_reset_reset_bridge_in_reset.reset
		.fpga_only_master_master_address                        (fpga_only_master_master_address),                                //                          fpga_only_master_master.address
		.fpga_only_master_master_waitrequest                    (fpga_only_master_master_waitrequest),                            //                                                 .waitrequest
		.fpga_only_master_master_byteenable                     (fpga_only_master_master_byteenable),                             //                                                 .byteenable
		.fpga_only_master_master_read                           (fpga_only_master_master_read),                                   //                                                 .read
		.fpga_only_master_master_readdata                       (fpga_only_master_master_readdata),                               //                                                 .readdata
		.fpga_only_master_master_readdatavalid                  (fpga_only_master_master_readdatavalid),                          //                                                 .readdatavalid
		.fpga_only_master_master_write                          (fpga_only_master_master_write),                                  //                                                 .write
		.fpga_only_master_master_writedata                      (fpga_only_master_master_writedata),                              //                                                 .writedata
		.mm_bridge_lw_axi_m0_address                            (mm_bridge_lw_axi_m0_address),                                    //                              mm_bridge_lw_axi_m0.address
		.mm_bridge_lw_axi_m0_waitrequest                        (mm_bridge_lw_axi_m0_waitrequest),                                //                                                 .waitrequest
		.mm_bridge_lw_axi_m0_burstcount                         (mm_bridge_lw_axi_m0_burstcount),                                 //                                                 .burstcount
		.mm_bridge_lw_axi_m0_byteenable                         (mm_bridge_lw_axi_m0_byteenable),                                 //                                                 .byteenable
		.mm_bridge_lw_axi_m0_read                               (mm_bridge_lw_axi_m0_read),                                       //                                                 .read
		.mm_bridge_lw_axi_m0_readdata                           (mm_bridge_lw_axi_m0_readdata),                                   //                                                 .readdata
		.mm_bridge_lw_axi_m0_readdatavalid                      (mm_bridge_lw_axi_m0_readdatavalid),                              //                                                 .readdatavalid
		.mm_bridge_lw_axi_m0_write                              (mm_bridge_lw_axi_m0_write),                                      //                                                 .write
		.mm_bridge_lw_axi_m0_writedata                          (mm_bridge_lw_axi_m0_writedata),                                  //                                                 .writedata
		.mm_bridge_lw_axi_m0_debugaccess                        (mm_bridge_lw_axi_m0_debugaccess),                                //                                                 .debugaccess
		.button_pio_s1_address                                  (mm_interconnect_3_button_pio_s1_address),                        //                                    button_pio_s1.address
		.button_pio_s1_write                                    (mm_interconnect_3_button_pio_s1_write),                          //                                                 .write
		.button_pio_s1_readdata                                 (mm_interconnect_3_button_pio_s1_readdata),                       //                                                 .readdata
		.button_pio_s1_writedata                                (mm_interconnect_3_button_pio_s1_writedata),                      //                                                 .writedata
		.button_pio_s1_chipselect                               (mm_interconnect_3_button_pio_s1_chipselect),                     //                                                 .chipselect
		.cnn_top_0_hps2cnn_avs_address                          (mm_interconnect_3_cnn_top_0_hps2cnn_avs_address),                //                            cnn_top_0_hps2cnn_avs.address
		.cnn_top_0_hps2cnn_avs_write                            (mm_interconnect_3_cnn_top_0_hps2cnn_avs_write),                  //                                                 .write
		.cnn_top_0_hps2cnn_avs_read                             (mm_interconnect_3_cnn_top_0_hps2cnn_avs_read),                   //                                                 .read
		.cnn_top_0_hps2cnn_avs_readdata                         (mm_interconnect_3_cnn_top_0_hps2cnn_avs_readdata),               //                                                 .readdata
		.cnn_top_0_hps2cnn_avs_writedata                        (mm_interconnect_3_cnn_top_0_hps2cnn_avs_writedata),              //                                                 .writedata
		.cnn_top_0_hps2cnn_avs_waitrequest                      (mm_interconnect_3_cnn_top_0_hps2cnn_avs_waitrequest),            //                                                 .waitrequest
		.ddr3_vga_0_cfg_bus_address                             (mm_interconnect_3_ddr3_vga_0_cfg_bus_address),                   //                               ddr3_vga_0_cfg_bus.address
		.ddr3_vga_0_cfg_bus_write                               (mm_interconnect_3_ddr3_vga_0_cfg_bus_write),                     //                                                 .write
		.ddr3_vga_0_cfg_bus_read                                (mm_interconnect_3_ddr3_vga_0_cfg_bus_read),                      //                                                 .read
		.ddr3_vga_0_cfg_bus_readdata                            (mm_interconnect_3_ddr3_vga_0_cfg_bus_readdata),                  //                                                 .readdata
		.ddr3_vga_0_cfg_bus_writedata                           (mm_interconnect_3_ddr3_vga_0_cfg_bus_writedata),                 //                                                 .writedata
		.dipsw_pio_s1_address                                   (mm_interconnect_3_dipsw_pio_s1_address),                         //                                     dipsw_pio_s1.address
		.dipsw_pio_s1_write                                     (mm_interconnect_3_dipsw_pio_s1_write),                           //                                                 .write
		.dipsw_pio_s1_readdata                                  (mm_interconnect_3_dipsw_pio_s1_readdata),                        //                                                 .readdata
		.dipsw_pio_s1_writedata                                 (mm_interconnect_3_dipsw_pio_s1_writedata),                       //                                                 .writedata
		.dipsw_pio_s1_chipselect                                (mm_interconnect_3_dipsw_pio_s1_chipselect),                      //                                                 .chipselect
		.dvp_ddr3_0_cfg_bus_address                             (mm_interconnect_3_dvp_ddr3_0_cfg_bus_address),                   //                               dvp_ddr3_0_cfg_bus.address
		.dvp_ddr3_0_cfg_bus_write                               (mm_interconnect_3_dvp_ddr3_0_cfg_bus_write),                     //                                                 .write
		.dvp_ddr3_0_cfg_bus_read                                (mm_interconnect_3_dvp_ddr3_0_cfg_bus_read),                      //                                                 .read
		.dvp_ddr3_0_cfg_bus_readdata                            (mm_interconnect_3_dvp_ddr3_0_cfg_bus_readdata),                  //                                                 .readdata
		.dvp_ddr3_0_cfg_bus_writedata                           (mm_interconnect_3_dvp_ddr3_0_cfg_bus_writedata),                 //                                                 .writedata
		.led_pio_s1_address                                     (mm_interconnect_3_led_pio_s1_address),                           //                                       led_pio_s1.address
		.led_pio_s1_write                                       (mm_interconnect_3_led_pio_s1_write),                             //                                                 .write
		.led_pio_s1_readdata                                    (mm_interconnect_3_led_pio_s1_readdata),                          //                                                 .readdata
		.led_pio_s1_writedata                                   (mm_interconnect_3_led_pio_s1_writedata),                         //                                                 .writedata
		.led_pio_s1_chipselect                                  (mm_interconnect_3_led_pio_s1_chipselect),                        //                                                 .chipselect
		.sld_hub_controller_system_0_s0_address                 (mm_interconnect_3_sld_hub_controller_system_0_s0_address),       //                   sld_hub_controller_system_0_s0.address
		.sld_hub_controller_system_0_s0_write                   (mm_interconnect_3_sld_hub_controller_system_0_s0_write),         //                                                 .write
		.sld_hub_controller_system_0_s0_read                    (mm_interconnect_3_sld_hub_controller_system_0_s0_read),          //                                                 .read
		.sld_hub_controller_system_0_s0_readdata                (mm_interconnect_3_sld_hub_controller_system_0_s0_readdata),      //                                                 .readdata
		.sld_hub_controller_system_0_s0_writedata               (mm_interconnect_3_sld_hub_controller_system_0_s0_writedata),     //                                                 .writedata
		.sld_hub_controller_system_0_s0_burstcount              (mm_interconnect_3_sld_hub_controller_system_0_s0_burstcount),    //                                                 .burstcount
		.sld_hub_controller_system_0_s0_byteenable              (mm_interconnect_3_sld_hub_controller_system_0_s0_byteenable),    //                                                 .byteenable
		.sld_hub_controller_system_0_s0_readdatavalid           (mm_interconnect_3_sld_hub_controller_system_0_s0_readdatavalid), //                                                 .readdatavalid
		.sld_hub_controller_system_0_s0_waitrequest             (mm_interconnect_3_sld_hub_controller_system_0_s0_waitrequest),   //                                                 .waitrequest
		.sld_hub_controller_system_0_s0_debugaccess             (mm_interconnect_3_sld_hub_controller_system_0_s0_debugaccess),   //                                                 .debugaccess
		.sysid_qsys_control_slave_address                       (mm_interconnect_3_sysid_qsys_control_slave_address),             //                         sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                      (mm_interconnect_3_sysid_qsys_control_slave_readdata),            //                                                 .readdata
		.vcam_0_cfg_bus_address                                 (mm_interconnect_3_vcam_0_cfg_bus_address),                       //                                   vcam_0_cfg_bus.address
		.vcam_0_cfg_bus_write                                   (mm_interconnect_3_vcam_0_cfg_bus_write),                         //                                                 .write
		.vcam_0_cfg_bus_read                                    (mm_interconnect_3_vcam_0_cfg_bus_read),                          //                                                 .read
		.vcam_0_cfg_bus_readdata                                (mm_interconnect_3_vcam_0_cfg_bus_readdata),                      //                                                 .readdata
		.vcam_0_cfg_bus_writedata                               (mm_interconnect_3_vcam_0_cfg_bus_writedata),                     //                                                 .writedata
		.vhdmi_0_s_avalon_mm_address                            (mm_interconnect_3_vhdmi_0_s_avalon_mm_address),                  //                              vhdmi_0_s_avalon_mm.address
		.vhdmi_0_s_avalon_mm_write                              (mm_interconnect_3_vhdmi_0_s_avalon_mm_write),                    //                                                 .write
		.vhdmi_0_s_avalon_mm_read                               (mm_interconnect_3_vhdmi_0_s_avalon_mm_read),                     //                                                 .read
		.vhdmi_0_s_avalon_mm_readdata                           (mm_interconnect_3_vhdmi_0_s_avalon_mm_readdata),                 //                                                 .readdata
		.vhdmi_0_s_avalon_mm_writedata                          (mm_interconnect_3_vhdmi_0_s_avalon_mm_writedata),                //                                                 .writedata
		.vhdmi_0_s_avalon_mm_chipselect                         (mm_interconnect_3_vhdmi_0_s_avalon_mm_chipselect)                //                                                 .chipselect
	);

	soc_system_mm_interconnect_4 mm_interconnect_4 (
		.hps_0_f2h_axi_slave_awid                                         (mm_interconnect_4_hps_0_f2h_axi_slave_awid),    //                                        hps_0_f2h_axi_slave.awid
		.hps_0_f2h_axi_slave_awaddr                                       (mm_interconnect_4_hps_0_f2h_axi_slave_awaddr),  //                                                           .awaddr
		.hps_0_f2h_axi_slave_awlen                                        (mm_interconnect_4_hps_0_f2h_axi_slave_awlen),   //                                                           .awlen
		.hps_0_f2h_axi_slave_awsize                                       (mm_interconnect_4_hps_0_f2h_axi_slave_awsize),  //                                                           .awsize
		.hps_0_f2h_axi_slave_awburst                                      (mm_interconnect_4_hps_0_f2h_axi_slave_awburst), //                                                           .awburst
		.hps_0_f2h_axi_slave_awlock                                       (mm_interconnect_4_hps_0_f2h_axi_slave_awlock),  //                                                           .awlock
		.hps_0_f2h_axi_slave_awcache                                      (mm_interconnect_4_hps_0_f2h_axi_slave_awcache), //                                                           .awcache
		.hps_0_f2h_axi_slave_awprot                                       (mm_interconnect_4_hps_0_f2h_axi_slave_awprot),  //                                                           .awprot
		.hps_0_f2h_axi_slave_awuser                                       (mm_interconnect_4_hps_0_f2h_axi_slave_awuser),  //                                                           .awuser
		.hps_0_f2h_axi_slave_awvalid                                      (mm_interconnect_4_hps_0_f2h_axi_slave_awvalid), //                                                           .awvalid
		.hps_0_f2h_axi_slave_awready                                      (mm_interconnect_4_hps_0_f2h_axi_slave_awready), //                                                           .awready
		.hps_0_f2h_axi_slave_wid                                          (mm_interconnect_4_hps_0_f2h_axi_slave_wid),     //                                                           .wid
		.hps_0_f2h_axi_slave_wdata                                        (mm_interconnect_4_hps_0_f2h_axi_slave_wdata),   //                                                           .wdata
		.hps_0_f2h_axi_slave_wstrb                                        (mm_interconnect_4_hps_0_f2h_axi_slave_wstrb),   //                                                           .wstrb
		.hps_0_f2h_axi_slave_wlast                                        (mm_interconnect_4_hps_0_f2h_axi_slave_wlast),   //                                                           .wlast
		.hps_0_f2h_axi_slave_wvalid                                       (mm_interconnect_4_hps_0_f2h_axi_slave_wvalid),  //                                                           .wvalid
		.hps_0_f2h_axi_slave_wready                                       (mm_interconnect_4_hps_0_f2h_axi_slave_wready),  //                                                           .wready
		.hps_0_f2h_axi_slave_bid                                          (mm_interconnect_4_hps_0_f2h_axi_slave_bid),     //                                                           .bid
		.hps_0_f2h_axi_slave_bresp                                        (mm_interconnect_4_hps_0_f2h_axi_slave_bresp),   //                                                           .bresp
		.hps_0_f2h_axi_slave_bvalid                                       (mm_interconnect_4_hps_0_f2h_axi_slave_bvalid),  //                                                           .bvalid
		.hps_0_f2h_axi_slave_bready                                       (mm_interconnect_4_hps_0_f2h_axi_slave_bready),  //                                                           .bready
		.hps_0_f2h_axi_slave_arid                                         (mm_interconnect_4_hps_0_f2h_axi_slave_arid),    //                                                           .arid
		.hps_0_f2h_axi_slave_araddr                                       (mm_interconnect_4_hps_0_f2h_axi_slave_araddr),  //                                                           .araddr
		.hps_0_f2h_axi_slave_arlen                                        (mm_interconnect_4_hps_0_f2h_axi_slave_arlen),   //                                                           .arlen
		.hps_0_f2h_axi_slave_arsize                                       (mm_interconnect_4_hps_0_f2h_axi_slave_arsize),  //                                                           .arsize
		.hps_0_f2h_axi_slave_arburst                                      (mm_interconnect_4_hps_0_f2h_axi_slave_arburst), //                                                           .arburst
		.hps_0_f2h_axi_slave_arlock                                       (mm_interconnect_4_hps_0_f2h_axi_slave_arlock),  //                                                           .arlock
		.hps_0_f2h_axi_slave_arcache                                      (mm_interconnect_4_hps_0_f2h_axi_slave_arcache), //                                                           .arcache
		.hps_0_f2h_axi_slave_arprot                                       (mm_interconnect_4_hps_0_f2h_axi_slave_arprot),  //                                                           .arprot
		.hps_0_f2h_axi_slave_aruser                                       (mm_interconnect_4_hps_0_f2h_axi_slave_aruser),  //                                                           .aruser
		.hps_0_f2h_axi_slave_arvalid                                      (mm_interconnect_4_hps_0_f2h_axi_slave_arvalid), //                                                           .arvalid
		.hps_0_f2h_axi_slave_arready                                      (mm_interconnect_4_hps_0_f2h_axi_slave_arready), //                                                           .arready
		.hps_0_f2h_axi_slave_rid                                          (mm_interconnect_4_hps_0_f2h_axi_slave_rid),     //                                                           .rid
		.hps_0_f2h_axi_slave_rdata                                        (mm_interconnect_4_hps_0_f2h_axi_slave_rdata),   //                                                           .rdata
		.hps_0_f2h_axi_slave_rresp                                        (mm_interconnect_4_hps_0_f2h_axi_slave_rresp),   //                                                           .rresp
		.hps_0_f2h_axi_slave_rlast                                        (mm_interconnect_4_hps_0_f2h_axi_slave_rlast),   //                                                           .rlast
		.hps_0_f2h_axi_slave_rvalid                                       (mm_interconnect_4_hps_0_f2h_axi_slave_rvalid),  //                                                           .rvalid
		.hps_0_f2h_axi_slave_rready                                       (mm_interconnect_4_hps_0_f2h_axi_slave_rready),  //                                                           .rready
		.clk_50_clk_clk                                                   (clk_50_clk),                                    //                                                 clk_50_clk.clk
		.hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),            // hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset.reset
		.hps_only_master_clk_reset_reset_bridge_in_reset_reset            (rst_controller_reset_out_reset),                //            hps_only_master_clk_reset_reset_bridge_in_reset.reset
		.mm_bridge_axi_reset_reset_bridge_in_reset_reset                  (rst_controller_reset_out_reset),                //                  mm_bridge_axi_reset_reset_bridge_in_reset.reset
		.hps_only_master_master_address                                   (hps_only_master_master_address),                //                                     hps_only_master_master.address
		.hps_only_master_master_waitrequest                               (hps_only_master_master_waitrequest),            //                                                           .waitrequest
		.hps_only_master_master_byteenable                                (hps_only_master_master_byteenable),             //                                                           .byteenable
		.hps_only_master_master_read                                      (hps_only_master_master_read),                   //                                                           .read
		.hps_only_master_master_readdata                                  (hps_only_master_master_readdata),               //                                                           .readdata
		.hps_only_master_master_readdatavalid                             (hps_only_master_master_readdatavalid),          //                                                           .readdatavalid
		.hps_only_master_master_write                                     (hps_only_master_master_write),                  //                                                           .write
		.hps_only_master_master_writedata                                 (hps_only_master_master_writedata),              //                                                           .writedata
		.mm_bridge_axi_m0_address                                         (mm_bridge_axi_m0_address),                      //                                           mm_bridge_axi_m0.address
		.mm_bridge_axi_m0_waitrequest                                     (mm_bridge_axi_m0_waitrequest),                  //                                                           .waitrequest
		.mm_bridge_axi_m0_burstcount                                      (mm_bridge_axi_m0_burstcount),                   //                                                           .burstcount
		.mm_bridge_axi_m0_byteenable                                      (mm_bridge_axi_m0_byteenable),                   //                                                           .byteenable
		.mm_bridge_axi_m0_read                                            (mm_bridge_axi_m0_read),                         //                                                           .read
		.mm_bridge_axi_m0_readdata                                        (mm_bridge_axi_m0_readdata),                     //                                                           .readdata
		.mm_bridge_axi_m0_readdatavalid                                   (mm_bridge_axi_m0_readdatavalid),                //                                                           .readdatavalid
		.mm_bridge_axi_m0_write                                           (mm_bridge_axi_m0_write),                        //                                                           .write
		.mm_bridge_axi_m0_writedata                                       (mm_bridge_axi_m0_writedata),                    //                                                           .writedata
		.mm_bridge_axi_m0_debugaccess                                     (mm_bridge_axi_m0_debugaccess)                   //                                                           .debugaccess
	);

	soc_system_mm_interconnect_5 mm_interconnect_5 (
		.clk_50_clk_clk                                                          (clk_50_clk),                                            //                                                        clk_50_clk.clk
		.clk_cnn_clk_clk                                                         (clk_cnn_clk),                                           //                                                       clk_cnn_clk.clk
		.f2sdram_only_master_clk_reset_reset_bridge_in_reset_reset               (rst_controller_reset_out_reset),                        //               f2sdram_only_master_clk_reset_reset_bridge_in_reset.reset
		.f2sdram_only_master_master_translator_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                        // f2sdram_only_master_master_translator_reset_reset_bridge_in_reset.reset
		.hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset      (rst_controller_003_reset_out_reset),                    //      hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset.reset
		.mm_bridge_sdram0_reset_reset_bridge_in_reset_reset                      (rst_controller_001_reset_out_reset),                    //                      mm_bridge_sdram0_reset_reset_bridge_in_reset.reset
		.f2sdram_only_master_master_address                                      (f2sdram_only_master_master_address),                    //                                        f2sdram_only_master_master.address
		.f2sdram_only_master_master_waitrequest                                  (f2sdram_only_master_master_waitrequest),                //                                                                  .waitrequest
		.f2sdram_only_master_master_byteenable                                   (f2sdram_only_master_master_byteenable),                 //                                                                  .byteenable
		.f2sdram_only_master_master_read                                         (f2sdram_only_master_master_read),                       //                                                                  .read
		.f2sdram_only_master_master_readdata                                     (f2sdram_only_master_master_readdata),                   //                                                                  .readdata
		.f2sdram_only_master_master_readdatavalid                                (f2sdram_only_master_master_readdatavalid),              //                                                                  .readdatavalid
		.f2sdram_only_master_master_write                                        (f2sdram_only_master_master_write),                      //                                                                  .write
		.f2sdram_only_master_master_writedata                                    (f2sdram_only_master_master_writedata),                  //                                                                  .writedata
		.mm_bridge_sdram0_m0_address                                             (mm_bridge_sdram0_m0_address),                           //                                               mm_bridge_sdram0_m0.address
		.mm_bridge_sdram0_m0_waitrequest                                         (mm_bridge_sdram0_m0_waitrequest),                       //                                                                  .waitrequest
		.mm_bridge_sdram0_m0_burstcount                                          (mm_bridge_sdram0_m0_burstcount),                        //                                                                  .burstcount
		.mm_bridge_sdram0_m0_byteenable                                          (mm_bridge_sdram0_m0_byteenable),                        //                                                                  .byteenable
		.mm_bridge_sdram0_m0_read                                                (mm_bridge_sdram0_m0_read),                              //                                                                  .read
		.mm_bridge_sdram0_m0_readdata                                            (mm_bridge_sdram0_m0_readdata),                          //                                                                  .readdata
		.mm_bridge_sdram0_m0_readdatavalid                                       (mm_bridge_sdram0_m0_readdatavalid),                     //                                                                  .readdatavalid
		.mm_bridge_sdram0_m0_write                                               (mm_bridge_sdram0_m0_write),                             //                                                                  .write
		.mm_bridge_sdram0_m0_writedata                                           (mm_bridge_sdram0_m0_writedata),                         //                                                                  .writedata
		.mm_bridge_sdram0_m0_debugaccess                                         (mm_bridge_sdram0_m0_debugaccess),                       //                                                                  .debugaccess
		.hps_0_f2h_sdram0_data_address                                           (mm_interconnect_5_hps_0_f2h_sdram0_data_address),       //                                             hps_0_f2h_sdram0_data.address
		.hps_0_f2h_sdram0_data_write                                             (mm_interconnect_5_hps_0_f2h_sdram0_data_write),         //                                                                  .write
		.hps_0_f2h_sdram0_data_read                                              (mm_interconnect_5_hps_0_f2h_sdram0_data_read),          //                                                                  .read
		.hps_0_f2h_sdram0_data_readdata                                          (mm_interconnect_5_hps_0_f2h_sdram0_data_readdata),      //                                                                  .readdata
		.hps_0_f2h_sdram0_data_writedata                                         (mm_interconnect_5_hps_0_f2h_sdram0_data_writedata),     //                                                                  .writedata
		.hps_0_f2h_sdram0_data_burstcount                                        (mm_interconnect_5_hps_0_f2h_sdram0_data_burstcount),    //                                                                  .burstcount
		.hps_0_f2h_sdram0_data_byteenable                                        (mm_interconnect_5_hps_0_f2h_sdram0_data_byteenable),    //                                                                  .byteenable
		.hps_0_f2h_sdram0_data_readdatavalid                                     (mm_interconnect_5_hps_0_f2h_sdram0_data_readdatavalid), //                                                                  .readdatavalid
		.hps_0_f2h_sdram0_data_waitrequest                                       (mm_interconnect_5_hps_0_f2h_sdram0_data_waitrequest)    //                                                                  .waitrequest
	);

	soc_system_irq_mapper irq_mapper (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq0_irq)  //    sender.irq
	);

	soc_system_irq_mapper irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_50_reset_n),              // reset_in0.reset
		.clk            (clk_50_clk),                     //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_cnn_reset_n),                 // reset_in0.reset
		.clk            (clk_cnn_clk),                        //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk            (clk_50_clk),                         //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk            (clk_cnn_clk),                        //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
